module Multiplexer_Hw( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [2:0]  io_5, // @[:@6.4]
  input         io_4_ready, // @[:@6.4]
  output        io_4_valid, // @[:@6.4]
  output [63:0] io_4_bits, // @[:@6.4]
  output        io_3_ready, // @[:@6.4]
  input         io_3_valid, // @[:@6.4]
  input  [63:0] io_3_bits, // @[:@6.4]
  output        io_2_ready, // @[:@6.4]
  input         io_2_valid, // @[:@6.4]
  input  [63:0] io_2_bits, // @[:@6.4]
  output        io_1_ready, // @[:@6.4]
  input         io_1_valid, // @[:@6.4]
  input  [63:0] io_1_bits, // @[:@6.4]
  output        io_0_ready, // @[:@6.4]
  input         io_0_valid, // @[:@6.4]
  input  [63:0] io_0_bits // @[:@6.4]
);
  wire [1:0] config$; // @[Multiplexer.scala 84:20:@8.4 Multiplexer.scala 85:10:@9.4]
  wire  _T_83; // @[Multiplexer.scala 105:17:@16.4]
  wire [63:0] _GEN_0; // @[Multiplexer.scala 105:30:@17.4]
  wire  _GEN_1; // @[Multiplexer.scala 105:30:@17.4]
  wire  _T_85; // @[Multiplexer.scala 105:17:@22.4]
  wire [63:0] _GEN_3; // @[Multiplexer.scala 105:30:@23.4]
  wire  _GEN_4; // @[Multiplexer.scala 105:30:@23.4]
  wire  _T_87; // @[Multiplexer.scala 105:17:@28.4]
  wire [63:0] _GEN_6; // @[Multiplexer.scala 105:30:@29.4]
  wire  _GEN_7; // @[Multiplexer.scala 105:30:@29.4]
  wire  _T_89; // @[Multiplexer.scala 105:17:@34.4]
  assign config$ = io_5[1:0]; // @[Multiplexer.scala 84:20:@8.4 Multiplexer.scala 85:10:@9.4]
  assign _T_83 = config$ == 2'h2; // @[Multiplexer.scala 105:17:@16.4]
  assign _GEN_0 = _T_83 ? io_2_bits : 64'h0; // @[Multiplexer.scala 105:30:@17.4]
  assign _GEN_1 = _T_83 ? io_2_valid : 1'h0; // @[Multiplexer.scala 105:30:@17.4]
  assign _T_85 = config$ == 2'h1; // @[Multiplexer.scala 105:17:@22.4]
  assign _GEN_3 = _T_85 ? io_1_bits : _GEN_0; // @[Multiplexer.scala 105:30:@23.4]
  assign _GEN_4 = _T_85 ? io_1_valid : _GEN_1; // @[Multiplexer.scala 105:30:@23.4]
  assign _T_87 = config$ == 2'h3; // @[Multiplexer.scala 105:17:@28.4]
  assign _GEN_6 = _T_87 ? io_3_bits : _GEN_3; // @[Multiplexer.scala 105:30:@29.4]
  assign _GEN_7 = _T_87 ? io_3_valid : _GEN_4; // @[Multiplexer.scala 105:30:@29.4]
  assign _T_89 = config$ == 2'h0; // @[Multiplexer.scala 105:17:@34.4]
  assign io_4_valid = _T_89 ? io_0_valid : _GEN_7; // @[Multiplexer.scala 91:28:@11.4 Multiplexer.scala 106:24:@19.6 Multiplexer.scala 106:24:@25.6 Multiplexer.scala 106:24:@31.6 Multiplexer.scala 106:24:@37.6]
  assign io_4_bits = _T_89 ? io_0_bits : _GEN_6; // @[Multiplexer.scala 91:13:@10.4 Multiplexer.scala 106:24:@18.6 Multiplexer.scala 106:24:@24.6 Multiplexer.scala 106:24:@30.6 Multiplexer.scala 106:24:@36.6]
  assign io_3_ready = _T_87 ? io_4_ready : 1'h0; // @[Multiplexer.scala 93:53:@15.4 Multiplexer.scala 106:24:@32.6]
  assign io_2_ready = _T_83 ? io_4_ready : 1'h0; // @[Multiplexer.scala 93:53:@14.4 Multiplexer.scala 106:24:@20.6]
  assign io_1_ready = _T_85 ? io_4_ready : 1'h0; // @[Multiplexer.scala 93:53:@13.4 Multiplexer.scala 106:24:@26.6]
  assign io_0_ready = _T_89 ? io_4_ready : 1'h0; // @[Multiplexer.scala 93:53:@12.4 Multiplexer.scala 106:24:@38.6]
endmodule
