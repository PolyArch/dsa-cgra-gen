module Delay_Pipe_Hw( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [2:0]  io_2, // @[:@6.4]
  output [31:0] io_1, // @[:@6.4]
  input  [31:0] io_0 // @[:@6.4]
);
  reg [2:0] head; // @[Delay_Pipe.scala 45:21:@8.4]
  reg [31:0] _RAND_0;
  reg [2:0] tail; // @[Delay_Pipe.scala 46:21:@9.4]
  reg [31:0] _RAND_1;
  reg [2:0] delay; // @[Delay_Pipe.scala 47:23:@10.4]
  reg [31:0] _RAND_2;
  reg [31:0] fifo_0; // @[Delay_Pipe.scala 50:21:@18.4]
  reg [31:0] _RAND_3;
  reg [31:0] fifo_1; // @[Delay_Pipe.scala 50:21:@18.4]
  reg [31:0] _RAND_4;
  reg [31:0] fifo_2; // @[Delay_Pipe.scala 50:21:@18.4]
  reg [31:0] _RAND_5;
  reg [31:0] fifo_3; // @[Delay_Pipe.scala 50:21:@18.4]
  reg [31:0] _RAND_6;
  reg [31:0] fifo_4; // @[Delay_Pipe.scala 50:21:@18.4]
  reg [31:0] _RAND_7;
  reg [31:0] fifo_5; // @[Delay_Pipe.scala 50:21:@18.4]
  reg [31:0] _RAND_8;
  wire [31:0] _GEN_1; // @[Delay_Pipe.scala 53:12:@19.4]
  wire [31:0] _GEN_2; // @[Delay_Pipe.scala 53:12:@19.4]
  wire [31:0] _GEN_3; // @[Delay_Pipe.scala 53:12:@19.4]
  wire [31:0] _GEN_4; // @[Delay_Pipe.scala 53:12:@19.4]
  wire [31:0] _GEN_6; // @[Delay_Pipe.scala 54:14:@20.4]
  wire [31:0] _GEN_7; // @[Delay_Pipe.scala 54:14:@20.4]
  wire [31:0] _GEN_8; // @[Delay_Pipe.scala 54:14:@20.4]
  wire [31:0] _GEN_9; // @[Delay_Pipe.scala 54:14:@20.4]
  wire [31:0] _GEN_10; // @[Delay_Pipe.scala 54:14:@20.4]
  wire [31:0] _GEN_11; // @[Delay_Pipe.scala 54:14:@20.4]
  wire [3:0] _T_83; // @[Delay_Pipe.scala 55:16:@21.4]
  wire [2:0] _T_84; // @[Delay_Pipe.scala 55:16:@22.4]
  wire [3:0] _T_86; // @[Delay_Pipe.scala 56:16:@24.4]
  wire [2:0] _T_87; // @[Delay_Pipe.scala 56:16:@25.4]
  wire  _T_88; // @[Delay_Pipe.scala 59:15:@27.4]
  wire [31:0] _GEN_12; // @[Delay_Pipe.scala 59:32:@28.4]
  wire [31:0] _GEN_13; // @[Delay_Pipe.scala 59:32:@28.4]
  wire [31:0] _GEN_14; // @[Delay_Pipe.scala 59:32:@28.4]
  wire [31:0] _GEN_15; // @[Delay_Pipe.scala 59:32:@28.4]
  wire [31:0] _GEN_16; // @[Delay_Pipe.scala 59:32:@28.4]
  wire [31:0] _GEN_17; // @[Delay_Pipe.scala 59:32:@28.4]
  wire [2:0] _GEN_18; // @[Delay_Pipe.scala 59:32:@28.4]
  wire [2:0] _GEN_19; // @[Delay_Pipe.scala 59:32:@28.4]
  assign _GEN_1 = 3'h1 == head ? fifo_1 : fifo_0; // @[Delay_Pipe.scala 53:12:@19.4]
  assign _GEN_2 = 3'h2 == head ? fifo_2 : _GEN_1; // @[Delay_Pipe.scala 53:12:@19.4]
  assign _GEN_3 = 3'h3 == head ? fifo_3 : _GEN_2; // @[Delay_Pipe.scala 53:12:@19.4]
  assign _GEN_4 = 3'h4 == head ? fifo_4 : _GEN_3; // @[Delay_Pipe.scala 53:12:@19.4]
  assign _GEN_6 = 3'h0 == tail ? io_0 : fifo_0; // @[Delay_Pipe.scala 54:14:@20.4]
  assign _GEN_7 = 3'h1 == tail ? io_0 : fifo_1; // @[Delay_Pipe.scala 54:14:@20.4]
  assign _GEN_8 = 3'h2 == tail ? io_0 : fifo_2; // @[Delay_Pipe.scala 54:14:@20.4]
  assign _GEN_9 = 3'h3 == tail ? io_0 : fifo_3; // @[Delay_Pipe.scala 54:14:@20.4]
  assign _GEN_10 = 3'h4 == tail ? io_0 : fifo_4; // @[Delay_Pipe.scala 54:14:@20.4]
  assign _GEN_11 = 3'h5 == tail ? io_0 : fifo_5; // @[Delay_Pipe.scala 54:14:@20.4]
  assign _T_83 = head + 3'h1; // @[Delay_Pipe.scala 55:16:@21.4]
  assign _T_84 = head + 3'h1; // @[Delay_Pipe.scala 55:16:@22.4]
  assign _T_86 = tail + 3'h1; // @[Delay_Pipe.scala 56:16:@24.4]
  assign _T_87 = tail + 3'h1; // @[Delay_Pipe.scala 56:16:@25.4]
  assign _T_88 = delay != io_2; // @[Delay_Pipe.scala 59:15:@27.4]
  assign _GEN_12 = _T_88 ? 32'h0 : _GEN_6; // @[Delay_Pipe.scala 59:32:@28.4]
  assign _GEN_13 = _T_88 ? 32'h0 : _GEN_7; // @[Delay_Pipe.scala 59:32:@28.4]
  assign _GEN_14 = _T_88 ? 32'h0 : _GEN_8; // @[Delay_Pipe.scala 59:32:@28.4]
  assign _GEN_15 = _T_88 ? 32'h0 : _GEN_9; // @[Delay_Pipe.scala 59:32:@28.4]
  assign _GEN_16 = _T_88 ? 32'h0 : _GEN_10; // @[Delay_Pipe.scala 59:32:@28.4]
  assign _GEN_17 = _T_88 ? 32'h0 : _GEN_11; // @[Delay_Pipe.scala 59:32:@28.4]
  assign _GEN_18 = _T_88 ? io_2 : _T_87; // @[Delay_Pipe.scala 59:32:@28.4]
  assign _GEN_19 = _T_88 ? io_2 : delay; // @[Delay_Pipe.scala 59:32:@28.4]
  assign io_1 = 3'h5 == head ? fifo_5 : _GEN_4; // @[Delay_Pipe.scala 53:12:@19.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  delay = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  fifo_0 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  fifo_1 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  fifo_2 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fifo_3 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  fifo_4 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  fifo_5 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      head <= 3'h0;
    end else begin
      head <= _T_84;
    end
    if (reset) begin
      tail <= 3'h0;
    end else begin
      if (_T_88) begin
        tail <= io_2;
      end else begin
        tail <= _T_87;
      end
    end
    if (reset) begin
      delay <= 3'h0;
    end else begin
      if (_T_88) begin
        delay <= io_2;
      end
    end
    if (reset) begin
      fifo_0 <= 32'h0;
    end else begin
      if (_T_88) begin
        fifo_0 <= 32'h0;
      end else begin
        if (3'h0 == tail) begin
          fifo_0 <= io_0;
        end
      end
    end
    if (reset) begin
      fifo_1 <= 32'h0;
    end else begin
      if (_T_88) begin
        fifo_1 <= 32'h0;
      end else begin
        if (3'h1 == tail) begin
          fifo_1 <= io_0;
        end
      end
    end
    if (reset) begin
      fifo_2 <= 32'h0;
    end else begin
      if (_T_88) begin
        fifo_2 <= 32'h0;
      end else begin
        if (3'h2 == tail) begin
          fifo_2 <= io_0;
        end
      end
    end
    if (reset) begin
      fifo_3 <= 32'h0;
    end else begin
      if (_T_88) begin
        fifo_3 <= 32'h0;
      end else begin
        if (3'h3 == tail) begin
          fifo_3 <= io_0;
        end
      end
    end
    if (reset) begin
      fifo_4 <= 32'h0;
    end else begin
      if (_T_88) begin
        fifo_4 <= 32'h0;
      end else begin
        if (3'h4 == tail) begin
          fifo_4 <= io_0;
        end
      end
    end
    if (reset) begin
      fifo_5 <= 32'h0;
    end else begin
      if (_T_88) begin
        fifo_5 <= 32'h0;
      end else begin
        if (3'h5 == tail) begin
          fifo_5 <= io_0;
        end
      end
    end
  end
endmodule
module Delay_Pipe_Hw_1( // @[:@39.2]
  input         clock, // @[:@40.4]
  input         reset, // @[:@41.4]
  input  [1:0]  io_2, // @[:@42.4]
  output [31:0] io_1, // @[:@42.4]
  input  [31:0] io_0 // @[:@42.4]
);
  reg [1:0] head; // @[Delay_Pipe.scala 45:21:@44.4]
  reg [31:0] _RAND_0;
  reg [1:0] tail; // @[Delay_Pipe.scala 46:21:@45.4]
  reg [31:0] _RAND_1;
  reg [1:0] delay; // @[Delay_Pipe.scala 47:23:@46.4]
  reg [31:0] _RAND_2;
  reg [31:0] fifo_0; // @[Delay_Pipe.scala 50:21:@51.4]
  reg [31:0] _RAND_3;
  reg [31:0] fifo_1; // @[Delay_Pipe.scala 50:21:@51.4]
  reg [31:0] _RAND_4;
  reg [31:0] fifo_2; // @[Delay_Pipe.scala 50:21:@51.4]
  reg [31:0] _RAND_5;
  wire [31:0] _GEN_1; // @[Delay_Pipe.scala 53:12:@52.4]
  wire [31:0] _GEN_3; // @[Delay_Pipe.scala 54:14:@53.4]
  wire [31:0] _GEN_4; // @[Delay_Pipe.scala 54:14:@53.4]
  wire [31:0] _GEN_5; // @[Delay_Pipe.scala 54:14:@53.4]
  wire [2:0] _T_62; // @[Delay_Pipe.scala 55:16:@54.4]
  wire [1:0] _T_63; // @[Delay_Pipe.scala 55:16:@55.4]
  wire [2:0] _T_65; // @[Delay_Pipe.scala 56:16:@57.4]
  wire [1:0] _T_66; // @[Delay_Pipe.scala 56:16:@58.4]
  wire  _T_67; // @[Delay_Pipe.scala 59:15:@60.4]
  wire [31:0] _GEN_6; // @[Delay_Pipe.scala 59:32:@61.4]
  wire [31:0] _GEN_7; // @[Delay_Pipe.scala 59:32:@61.4]
  wire [31:0] _GEN_8; // @[Delay_Pipe.scala 59:32:@61.4]
  wire [1:0] _GEN_9; // @[Delay_Pipe.scala 59:32:@61.4]
  wire [1:0] _GEN_10; // @[Delay_Pipe.scala 59:32:@61.4]
  assign _GEN_1 = 2'h1 == head ? fifo_1 : fifo_0; // @[Delay_Pipe.scala 53:12:@52.4]
  assign _GEN_3 = 2'h0 == tail ? io_0 : fifo_0; // @[Delay_Pipe.scala 54:14:@53.4]
  assign _GEN_4 = 2'h1 == tail ? io_0 : fifo_1; // @[Delay_Pipe.scala 54:14:@53.4]
  assign _GEN_5 = 2'h2 == tail ? io_0 : fifo_2; // @[Delay_Pipe.scala 54:14:@53.4]
  assign _T_62 = head + 2'h1; // @[Delay_Pipe.scala 55:16:@54.4]
  assign _T_63 = head + 2'h1; // @[Delay_Pipe.scala 55:16:@55.4]
  assign _T_65 = tail + 2'h1; // @[Delay_Pipe.scala 56:16:@57.4]
  assign _T_66 = tail + 2'h1; // @[Delay_Pipe.scala 56:16:@58.4]
  assign _T_67 = delay != io_2; // @[Delay_Pipe.scala 59:15:@60.4]
  assign _GEN_6 = _T_67 ? 32'h0 : _GEN_3; // @[Delay_Pipe.scala 59:32:@61.4]
  assign _GEN_7 = _T_67 ? 32'h0 : _GEN_4; // @[Delay_Pipe.scala 59:32:@61.4]
  assign _GEN_8 = _T_67 ? 32'h0 : _GEN_5; // @[Delay_Pipe.scala 59:32:@61.4]
  assign _GEN_9 = _T_67 ? io_2 : _T_66; // @[Delay_Pipe.scala 59:32:@61.4]
  assign _GEN_10 = _T_67 ? io_2 : delay; // @[Delay_Pipe.scala 59:32:@61.4]
  assign io_1 = 2'h2 == head ? fifo_2 : _GEN_1; // @[Delay_Pipe.scala 53:12:@52.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  delay = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  fifo_0 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  fifo_1 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  fifo_2 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      head <= 2'h0;
    end else begin
      head <= _T_63;
    end
    if (reset) begin
      tail <= 2'h0;
    end else begin
      if (_T_67) begin
        tail <= io_2;
      end else begin
        tail <= _T_66;
      end
    end
    if (reset) begin
      delay <= 2'h0;
    end else begin
      if (_T_67) begin
        delay <= io_2;
      end
    end
    if (reset) begin
      fifo_0 <= 32'h0;
    end else begin
      if (_T_67) begin
        fifo_0 <= 32'h0;
      end else begin
        if (2'h0 == tail) begin
          fifo_0 <= io_0;
        end
      end
    end
    if (reset) begin
      fifo_1 <= 32'h0;
    end else begin
      if (_T_67) begin
        fifo_1 <= 32'h0;
      end else begin
        if (2'h1 == tail) begin
          fifo_1 <= io_0;
        end
      end
    end
    if (reset) begin
      fifo_2 <= 32'h0;
    end else begin
      if (_T_67) begin
        fifo_2 <= 32'h0;
      end else begin
        if (2'h2 == tail) begin
          fifo_2 <= io_0;
        end
      end
    end
  end
endmodule
module Arithmetic_Logic_Unit_Hw( // @[:@99.2]
  input         clock, // @[:@100.4]
  input         reset, // @[:@101.4]
  input  [4:0]  io_4, // @[:@102.4]
  input  [31:0] io_3, // @[:@102.4]
  output [31:0] io_2, // @[:@102.4]
  input  [31:0] io_1, // @[:@102.4]
  input  [31:0] io_0 // @[:@102.4]
);
  wire  logical_operand0_unsigned; // @[Arithmetic_Logic_Unit.scala 91:58:@127.4]
  wire  logical_operand1_unsigned; // @[Arithmetic_Logic_Unit.scala 92:58:@128.4]
  wire  logical_operand2_unsigned; // @[Arithmetic_Logic_Unit.scala 93:58:@129.4]
  wire  _T_43; // @[Arithmetic_Logic_Unit.scala 96:49:@134.4]
  wire [31:0] _GEN_1; // @[Arithmetic_Logic_Unit.scala 96:65:@135.4]
  wire  _T_45; // @[Arithmetic_Logic_Unit.scala 97:49:@138.4]
  wire [32:0] _T_46; // @[Arithmetic_Logic_Unit.scala 97:103:@140.6]
  wire [31:0] _T_47; // @[Arithmetic_Logic_Unit.scala 97:103:@141.6]
  wire [31:0] _GEN_2; // @[Arithmetic_Logic_Unit.scala 97:65:@139.4]
  wire  _T_49; // @[Arithmetic_Logic_Unit.scala 98:49:@144.4]
  wire [32:0] _T_50; // @[Arithmetic_Logic_Unit.scala 98:103:@146.6]
  wire [32:0] _T_51; // @[Arithmetic_Logic_Unit.scala 98:103:@147.6]
  wire [31:0] _T_52; // @[Arithmetic_Logic_Unit.scala 98:103:@148.6]
  wire [31:0] _GEN_3; // @[Arithmetic_Logic_Unit.scala 98:65:@145.4]
  wire  _T_54; // @[Arithmetic_Logic_Unit.scala 99:49:@151.4]
  wire [18:0] _T_55; // @[Arithmetic_Logic_Unit.scala 99:123:@153.6]
  wire [524318:0] _GEN_37; // @[Arithmetic_Logic_Unit.scala 99:103:@154.6]
  wire [524318:0] _T_56; // @[Arithmetic_Logic_Unit.scala 99:103:@154.6]
  wire [524318:0] _GEN_4; // @[Arithmetic_Logic_Unit.scala 99:65:@152.4]
  wire  _T_58; // @[Arithmetic_Logic_Unit.scala 100:49:@157.4]
  wire [31:0] _T_59; // @[Arithmetic_Logic_Unit.scala 100:103:@159.6]
  wire [524318:0] _GEN_5; // @[Arithmetic_Logic_Unit.scala 100:65:@158.4]
  wire  _T_61; // @[Arithmetic_Logic_Unit.scala 101:48:@162.4]
  wire  _T_62; // @[Arithmetic_Logic_Unit.scala 101:101:@164.6]
  wire [524318:0] _GEN_6; // @[Arithmetic_Logic_Unit.scala 101:63:@163.4]
  wire  _T_64; // @[Arithmetic_Logic_Unit.scala 102:48:@167.4]
  wire  _T_65; // @[Arithmetic_Logic_Unit.scala 102:101:@169.6]
  wire [524318:0] _GEN_7; // @[Arithmetic_Logic_Unit.scala 102:63:@168.4]
  wire  _T_67; // @[Arithmetic_Logic_Unit.scala 103:49:@172.4]
  wire  _T_68; // @[Arithmetic_Logic_Unit.scala 103:103:@174.6]
  wire [524318:0] _GEN_8; // @[Arithmetic_Logic_Unit.scala 103:65:@173.4]
  wire  _T_70; // @[Arithmetic_Logic_Unit.scala 104:49:@177.4]
  wire  _T_71; // @[Arithmetic_Logic_Unit.scala 104:104:@179.6]
  wire [524318:0] _GEN_9; // @[Arithmetic_Logic_Unit.scala 104:66:@178.4]
  wire  _T_73; // @[Arithmetic_Logic_Unit.scala 105:49:@182.4]
  wire  _T_74; // @[Arithmetic_Logic_Unit.scala 105:103:@184.6]
  wire [524318:0] _GEN_10; // @[Arithmetic_Logic_Unit.scala 105:65:@183.4]
  wire  _T_76; // @[Arithmetic_Logic_Unit.scala 106:49:@187.4]
  wire  _T_77; // @[Arithmetic_Logic_Unit.scala 106:103:@189.6]
  wire [524318:0] _GEN_11; // @[Arithmetic_Logic_Unit.scala 106:65:@188.4]
  wire  _T_79; // @[Arithmetic_Logic_Unit.scala 107:50:@192.4]
  wire [31:0] _T_80; // @[Arithmetic_Logic_Unit.scala 107:105:@194.6]
  wire [524318:0] _GEN_12; // @[Arithmetic_Logic_Unit.scala 107:67:@193.4]
  wire  _T_82; // @[Arithmetic_Logic_Unit.scala 108:51:@197.4]
  wire [31:0] _T_84; // @[Arithmetic_Logic_Unit.scala 108:89:@200.6]
  wire [524318:0] _GEN_13; // @[Arithmetic_Logic_Unit.scala 108:69:@198.4]
  wire  _T_86; // @[Arithmetic_Logic_Unit.scala 109:49:@203.4]
  wire [31:0] _T_87; // @[Arithmetic_Logic_Unit.scala 109:103:@205.6]
  wire [524318:0] _GEN_14; // @[Arithmetic_Logic_Unit.scala 109:65:@204.4]
  wire  _T_89; // @[Arithmetic_Logic_Unit.scala 110:50:@208.4]
  wire [31:0] _T_91; // @[Arithmetic_Logic_Unit.scala 110:87:@211.6]
  wire [524318:0] _GEN_15; // @[Arithmetic_Logic_Unit.scala 110:67:@209.4]
  wire  _T_93; // @[Arithmetic_Logic_Unit.scala 111:50:@214.4]
  wire [31:0] _T_94; // @[Arithmetic_Logic_Unit.scala 111:105:@216.6]
  wire [524318:0] _GEN_16; // @[Arithmetic_Logic_Unit.scala 111:67:@215.4]
  wire  _T_96; // @[Arithmetic_Logic_Unit.scala 112:51:@219.4]
  wire [31:0] _T_98; // @[Arithmetic_Logic_Unit.scala 112:89:@222.6]
  wire [524318:0] _GEN_17; // @[Arithmetic_Logic_Unit.scala 112:69:@220.4]
  wire  _T_100; // @[Arithmetic_Logic_Unit.scala 113:50:@225.4]
  wire  _T_101; // @[Arithmetic_Logic_Unit.scala 113:113:@227.6]
  wire [524318:0] _GEN_18; // @[Arithmetic_Logic_Unit.scala 113:67:@226.4]
  wire  _T_103; // @[Arithmetic_Logic_Unit.scala 114:51:@230.4]
  wire  _T_106; // @[Arithmetic_Logic_Unit.scala 114:89:@233.6]
  wire [524318:0] _GEN_19; // @[Arithmetic_Logic_Unit.scala 114:69:@231.4]
  wire  _T_108; // @[Arithmetic_Logic_Unit.scala 115:49:@236.4]
  wire  _T_109; // @[Arithmetic_Logic_Unit.scala 115:111:@238.6]
  wire [524318:0] _GEN_20; // @[Arithmetic_Logic_Unit.scala 115:65:@237.4]
  wire  _T_111; // @[Arithmetic_Logic_Unit.scala 116:50:@241.4]
  wire  _T_114; // @[Arithmetic_Logic_Unit.scala 116:87:@244.6]
  wire [524318:0] _GEN_21; // @[Arithmetic_Logic_Unit.scala 116:67:@242.4]
  wire  _T_116; // @[Arithmetic_Logic_Unit.scala 117:50:@247.4]
  wire  _T_118; // @[Arithmetic_Logic_Unit.scala 117:87:@249.6]
  wire  _T_120; // @[Arithmetic_Logic_Unit.scala 117:116:@250.6]
  wire  _T_121; // @[Arithmetic_Logic_Unit.scala 117:114:@251.6]
  wire [524318:0] _GEN_22; // @[Arithmetic_Logic_Unit.scala 117:67:@248.4]
  wire  _T_123; // @[Arithmetic_Logic_Unit.scala 118:51:@254.4]
  wire  _T_130; // @[Arithmetic_Logic_Unit.scala 118:89:@259.6]
  wire [524318:0] _GEN_23; // @[Arithmetic_Logic_Unit.scala 118:69:@255.4]
  wire [5:0] _GEN_38; // @[Arithmetic_Logic_Unit.scala 119:48:@262.4]
  wire  _T_132; // @[Arithmetic_Logic_Unit.scala 119:48:@262.4]
  wire  _T_134; // @[Arithmetic_Logic_Unit.scala 119:100:@265.6]
  wire [524318:0] _GEN_24; // @[Arithmetic_Logic_Unit.scala 119:63:@263.4]
  wire  _T_136; // @[Arithmetic_Logic_Unit.scala 120:48:@268.4]
  wire [524287:0] _T_139; // @[Arithmetic_Logic_Unit.scala 122:53:@272.8]
  wire [524287:0] _GEN_40; // @[Arithmetic_Logic_Unit.scala 122:46:@273.8]
  wire [524287:0] _T_140; // @[Arithmetic_Logic_Unit.scala 122:46:@273.8]
  wire [524287:0] _T_144; // @[Arithmetic_Logic_Unit.scala 124:49:@279.8]
  wire [524287:0] _T_145; // @[Arithmetic_Logic_Unit.scala 124:46:@280.8]
  wire [524287:0] _GEN_25; // @[Arithmetic_Logic_Unit.scala 121:38:@270.6]
  wire [524318:0] _GEN_26; // @[Arithmetic_Logic_Unit.scala 120:63:@269.4]
  wire  _T_147; // @[Arithmetic_Logic_Unit.scala 127:48:@284.4]
  wire [524318:0] _GEN_27; // @[Arithmetic_Logic_Unit.scala 127:63:@285.4]
  wire  _T_154; // @[Arithmetic_Logic_Unit.scala 128:48:@292.4]
  wire [524318:0] _GEN_28; // @[Arithmetic_Logic_Unit.scala 128:63:@293.4]
  wire  _T_160; // @[Arithmetic_Logic_Unit.scala 129:49:@299.4]
  wire  _T_162; // @[Arithmetic_Logic_Unit.scala 130:30:@301.6]
  wire [15:0] _T_168; // @[Bitwise.scala 103:21:@308.8]
  wire [31:0] _T_169; // @[Bitwise.scala 103:31:@309.8]
  wire [15:0] _T_170; // @[Bitwise.scala 103:46:@310.8]
  wire [31:0] _GEN_47; // @[Bitwise.scala 103:65:@311.8]
  wire [31:0] _T_171; // @[Bitwise.scala 103:65:@311.8]
  wire [31:0] _T_173; // @[Bitwise.scala 103:75:@313.8]
  wire [31:0] _T_174; // @[Bitwise.scala 103:39:@314.8]
  wire [23:0] _T_178; // @[Bitwise.scala 103:21:@318.8]
  wire [31:0] _GEN_48; // @[Bitwise.scala 103:31:@319.8]
  wire [31:0] _T_179; // @[Bitwise.scala 103:31:@319.8]
  wire [23:0] _T_180; // @[Bitwise.scala 103:46:@320.8]
  wire [31:0] _GEN_49; // @[Bitwise.scala 103:65:@321.8]
  wire [31:0] _T_181; // @[Bitwise.scala 103:65:@321.8]
  wire [31:0] _T_183; // @[Bitwise.scala 103:75:@323.8]
  wire [31:0] _T_184; // @[Bitwise.scala 103:39:@324.8]
  wire [27:0] _T_188; // @[Bitwise.scala 103:21:@328.8]
  wire [31:0] _GEN_50; // @[Bitwise.scala 103:31:@329.8]
  wire [31:0] _T_189; // @[Bitwise.scala 103:31:@329.8]
  wire [27:0] _T_190; // @[Bitwise.scala 103:46:@330.8]
  wire [31:0] _GEN_51; // @[Bitwise.scala 103:65:@331.8]
  wire [31:0] _T_191; // @[Bitwise.scala 103:65:@331.8]
  wire [31:0] _T_193; // @[Bitwise.scala 103:75:@333.8]
  wire [31:0] _T_194; // @[Bitwise.scala 103:39:@334.8]
  wire [29:0] _T_198; // @[Bitwise.scala 103:21:@338.8]
  wire [31:0] _GEN_52; // @[Bitwise.scala 103:31:@339.8]
  wire [31:0] _T_199; // @[Bitwise.scala 103:31:@339.8]
  wire [29:0] _T_200; // @[Bitwise.scala 103:46:@340.8]
  wire [31:0] _GEN_53; // @[Bitwise.scala 103:65:@341.8]
  wire [31:0] _T_201; // @[Bitwise.scala 103:65:@341.8]
  wire [31:0] _T_203; // @[Bitwise.scala 103:75:@343.8]
  wire [31:0] _T_204; // @[Bitwise.scala 103:39:@344.8]
  wire [30:0] _T_208; // @[Bitwise.scala 103:21:@348.8]
  wire [31:0] _GEN_54; // @[Bitwise.scala 103:31:@349.8]
  wire [31:0] _T_209; // @[Bitwise.scala 103:31:@349.8]
  wire [30:0] _T_210; // @[Bitwise.scala 103:46:@350.8]
  wire [31:0] _GEN_55; // @[Bitwise.scala 103:65:@351.8]
  wire [31:0] _T_211; // @[Bitwise.scala 103:65:@351.8]
  wire [31:0] _T_213; // @[Bitwise.scala 103:75:@353.8]
  wire [31:0] _T_214; // @[Bitwise.scala 103:39:@354.8]
  wire  _T_215; // @[OneHot.scala 39:40:@355.8]
  wire  _T_216; // @[OneHot.scala 39:40:@356.8]
  wire  _T_217; // @[OneHot.scala 39:40:@357.8]
  wire  _T_218; // @[OneHot.scala 39:40:@358.8]
  wire  _T_219; // @[OneHot.scala 39:40:@359.8]
  wire  _T_220; // @[OneHot.scala 39:40:@360.8]
  wire  _T_221; // @[OneHot.scala 39:40:@361.8]
  wire  _T_222; // @[OneHot.scala 39:40:@362.8]
  wire  _T_223; // @[OneHot.scala 39:40:@363.8]
  wire  _T_224; // @[OneHot.scala 39:40:@364.8]
  wire  _T_225; // @[OneHot.scala 39:40:@365.8]
  wire  _T_226; // @[OneHot.scala 39:40:@366.8]
  wire  _T_227; // @[OneHot.scala 39:40:@367.8]
  wire  _T_228; // @[OneHot.scala 39:40:@368.8]
  wire  _T_229; // @[OneHot.scala 39:40:@369.8]
  wire  _T_230; // @[OneHot.scala 39:40:@370.8]
  wire  _T_231; // @[OneHot.scala 39:40:@371.8]
  wire  _T_232; // @[OneHot.scala 39:40:@372.8]
  wire  _T_233; // @[OneHot.scala 39:40:@373.8]
  wire  _T_234; // @[OneHot.scala 39:40:@374.8]
  wire  _T_235; // @[OneHot.scala 39:40:@375.8]
  wire  _T_236; // @[OneHot.scala 39:40:@376.8]
  wire  _T_237; // @[OneHot.scala 39:40:@377.8]
  wire  _T_238; // @[OneHot.scala 39:40:@378.8]
  wire  _T_239; // @[OneHot.scala 39:40:@379.8]
  wire  _T_240; // @[OneHot.scala 39:40:@380.8]
  wire  _T_241; // @[OneHot.scala 39:40:@381.8]
  wire  _T_242; // @[OneHot.scala 39:40:@382.8]
  wire  _T_243; // @[OneHot.scala 39:40:@383.8]
  wire  _T_244; // @[OneHot.scala 39:40:@384.8]
  wire  _T_245; // @[OneHot.scala 39:40:@385.8]
  wire [4:0] _T_279; // @[Mux.scala 31:69:@387.8]
  wire [4:0] _T_280; // @[Mux.scala 31:69:@388.8]
  wire [4:0] _T_281; // @[Mux.scala 31:69:@389.8]
  wire [4:0] _T_282; // @[Mux.scala 31:69:@390.8]
  wire [4:0] _T_283; // @[Mux.scala 31:69:@391.8]
  wire [4:0] _T_284; // @[Mux.scala 31:69:@392.8]
  wire [4:0] _T_285; // @[Mux.scala 31:69:@393.8]
  wire [4:0] _T_286; // @[Mux.scala 31:69:@394.8]
  wire [4:0] _T_287; // @[Mux.scala 31:69:@395.8]
  wire [4:0] _T_288; // @[Mux.scala 31:69:@396.8]
  wire [4:0] _T_289; // @[Mux.scala 31:69:@397.8]
  wire [4:0] _T_290; // @[Mux.scala 31:69:@398.8]
  wire [4:0] _T_291; // @[Mux.scala 31:69:@399.8]
  wire [4:0] _T_292; // @[Mux.scala 31:69:@400.8]
  wire [4:0] _T_293; // @[Mux.scala 31:69:@401.8]
  wire [4:0] _T_294; // @[Mux.scala 31:69:@402.8]
  wire [4:0] _T_295; // @[Mux.scala 31:69:@403.8]
  wire [4:0] _T_296; // @[Mux.scala 31:69:@404.8]
  wire [4:0] _T_297; // @[Mux.scala 31:69:@405.8]
  wire [4:0] _T_298; // @[Mux.scala 31:69:@406.8]
  wire [4:0] _T_299; // @[Mux.scala 31:69:@407.8]
  wire [4:0] _T_300; // @[Mux.scala 31:69:@408.8]
  wire [4:0] _T_301; // @[Mux.scala 31:69:@409.8]
  wire [4:0] _T_302; // @[Mux.scala 31:69:@410.8]
  wire [4:0] _T_303; // @[Mux.scala 31:69:@411.8]
  wire [4:0] _T_304; // @[Mux.scala 31:69:@412.8]
  wire [4:0] _T_305; // @[Mux.scala 31:69:@413.8]
  wire [4:0] _T_306; // @[Mux.scala 31:69:@414.8]
  wire [4:0] _T_307; // @[Mux.scala 31:69:@415.8]
  wire [4:0] _T_308; // @[Mux.scala 31:69:@416.8]
  wire [4:0] _T_309; // @[Mux.scala 31:69:@417.8]
  wire [5:0] _GEN_29; // @[Arithmetic_Logic_Unit.scala 130:38:@302.6]
  wire [524318:0] _GEN_30; // @[Arithmetic_Logic_Unit.scala 129:65:@300.4]
  wire  _T_311; // @[Arithmetic_Logic_Unit.scala 136:49:@421.4]
  wire  _T_315; // @[OneHot.scala 39:40:@428.8]
  wire  _T_316; // @[OneHot.scala 39:40:@429.8]
  wire  _T_317; // @[OneHot.scala 39:40:@430.8]
  wire  _T_318; // @[OneHot.scala 39:40:@431.8]
  wire  _T_319; // @[OneHot.scala 39:40:@432.8]
  wire  _T_320; // @[OneHot.scala 39:40:@433.8]
  wire  _T_321; // @[OneHot.scala 39:40:@434.8]
  wire  _T_322; // @[OneHot.scala 39:40:@435.8]
  wire  _T_323; // @[OneHot.scala 39:40:@436.8]
  wire  _T_324; // @[OneHot.scala 39:40:@437.8]
  wire  _T_325; // @[OneHot.scala 39:40:@438.8]
  wire  _T_326; // @[OneHot.scala 39:40:@439.8]
  wire  _T_327; // @[OneHot.scala 39:40:@440.8]
  wire  _T_328; // @[OneHot.scala 39:40:@441.8]
  wire  _T_329; // @[OneHot.scala 39:40:@442.8]
  wire  _T_330; // @[OneHot.scala 39:40:@443.8]
  wire  _T_331; // @[OneHot.scala 39:40:@444.8]
  wire  _T_332; // @[OneHot.scala 39:40:@445.8]
  wire  _T_333; // @[OneHot.scala 39:40:@446.8]
  wire  _T_334; // @[OneHot.scala 39:40:@447.8]
  wire  _T_335; // @[OneHot.scala 39:40:@448.8]
  wire  _T_336; // @[OneHot.scala 39:40:@449.8]
  wire  _T_337; // @[OneHot.scala 39:40:@450.8]
  wire  _T_338; // @[OneHot.scala 39:40:@451.8]
  wire  _T_339; // @[OneHot.scala 39:40:@452.8]
  wire  _T_340; // @[OneHot.scala 39:40:@453.8]
  wire  _T_341; // @[OneHot.scala 39:40:@454.8]
  wire  _T_342; // @[OneHot.scala 39:40:@455.8]
  wire  _T_343; // @[OneHot.scala 39:40:@456.8]
  wire  _T_344; // @[OneHot.scala 39:40:@457.8]
  wire  _T_345; // @[OneHot.scala 39:40:@458.8]
  wire [4:0] _T_379; // @[Mux.scala 31:69:@460.8]
  wire [4:0] _T_380; // @[Mux.scala 31:69:@461.8]
  wire [4:0] _T_381; // @[Mux.scala 31:69:@462.8]
  wire [4:0] _T_382; // @[Mux.scala 31:69:@463.8]
  wire [4:0] _T_383; // @[Mux.scala 31:69:@464.8]
  wire [4:0] _T_384; // @[Mux.scala 31:69:@465.8]
  wire [4:0] _T_385; // @[Mux.scala 31:69:@466.8]
  wire [4:0] _T_386; // @[Mux.scala 31:69:@467.8]
  wire [4:0] _T_387; // @[Mux.scala 31:69:@468.8]
  wire [4:0] _T_388; // @[Mux.scala 31:69:@469.8]
  wire [4:0] _T_389; // @[Mux.scala 31:69:@470.8]
  wire [4:0] _T_390; // @[Mux.scala 31:69:@471.8]
  wire [4:0] _T_391; // @[Mux.scala 31:69:@472.8]
  wire [4:0] _T_392; // @[Mux.scala 31:69:@473.8]
  wire [4:0] _T_393; // @[Mux.scala 31:69:@474.8]
  wire [4:0] _T_394; // @[Mux.scala 31:69:@475.8]
  wire [4:0] _T_395; // @[Mux.scala 31:69:@476.8]
  wire [4:0] _T_396; // @[Mux.scala 31:69:@477.8]
  wire [4:0] _T_397; // @[Mux.scala 31:69:@478.8]
  wire [4:0] _T_398; // @[Mux.scala 31:69:@479.8]
  wire [4:0] _T_399; // @[Mux.scala 31:69:@480.8]
  wire [4:0] _T_400; // @[Mux.scala 31:69:@481.8]
  wire [4:0] _T_401; // @[Mux.scala 31:69:@482.8]
  wire [4:0] _T_402; // @[Mux.scala 31:69:@483.8]
  wire [4:0] _T_403; // @[Mux.scala 31:69:@484.8]
  wire [4:0] _T_404; // @[Mux.scala 31:69:@485.8]
  wire [4:0] _T_405; // @[Mux.scala 31:69:@486.8]
  wire [4:0] _T_406; // @[Mux.scala 31:69:@487.8]
  wire [4:0] _T_407; // @[Mux.scala 31:69:@488.8]
  wire [4:0] _T_408; // @[Mux.scala 31:69:@489.8]
  wire [4:0] _T_409; // @[Mux.scala 31:69:@490.8]
  wire [5:0] _GEN_31; // @[Arithmetic_Logic_Unit.scala 137:39:@424.6]
  wire [524318:0] _GEN_32; // @[Arithmetic_Logic_Unit.scala 136:65:@422.4]
  wire  _T_411; // @[Arithmetic_Logic_Unit.scala 143:50:@494.4]
  wire [524318:0] _GEN_33; // @[Arithmetic_Logic_Unit.scala 143:67:@495.4]
  wire  _T_483; // @[Arithmetic_Logic_Unit.scala 171:58:@532.4]
  wire  _T_484; // @[Arithmetic_Logic_Unit.scala 171:58:@533.4]
  wire  _T_485; // @[Arithmetic_Logic_Unit.scala 171:58:@534.4]
  wire  _T_486; // @[Arithmetic_Logic_Unit.scala 171:58:@535.4]
  wire  _T_487; // @[Arithmetic_Logic_Unit.scala 171:58:@536.4]
  wire  _T_488; // @[Arithmetic_Logic_Unit.scala 171:58:@537.4]
  wire  _T_489; // @[Arithmetic_Logic_Unit.scala 171:58:@538.4]
  wire  _T_490; // @[Arithmetic_Logic_Unit.scala 171:58:@539.4]
  wire  _T_491; // @[Arithmetic_Logic_Unit.scala 171:58:@540.4]
  wire  _T_492; // @[Arithmetic_Logic_Unit.scala 171:58:@541.4]
  wire  _T_493; // @[Arithmetic_Logic_Unit.scala 171:58:@542.4]
  wire  _T_494; // @[Arithmetic_Logic_Unit.scala 171:58:@543.4]
  wire  _T_495; // @[Arithmetic_Logic_Unit.scala 171:58:@544.4]
  wire  _T_496; // @[Arithmetic_Logic_Unit.scala 171:58:@545.4]
  wire  _T_497; // @[Arithmetic_Logic_Unit.scala 171:58:@546.4]
  wire  _T_498; // @[Arithmetic_Logic_Unit.scala 171:58:@547.4]
  wire  _T_499; // @[Arithmetic_Logic_Unit.scala 171:58:@548.4]
  wire  _T_500; // @[Arithmetic_Logic_Unit.scala 171:58:@549.4]
  wire  _T_501; // @[Arithmetic_Logic_Unit.scala 171:58:@550.4]
  wire  _T_502; // @[Arithmetic_Logic_Unit.scala 171:58:@551.4]
  wire  _T_503; // @[Arithmetic_Logic_Unit.scala 171:58:@552.4]
  wire  _T_504; // @[Arithmetic_Logic_Unit.scala 171:58:@553.4]
  wire  _T_505; // @[Arithmetic_Logic_Unit.scala 171:58:@554.4]
  wire  _T_506; // @[Arithmetic_Logic_Unit.scala 171:58:@555.4]
  wire  _T_507; // @[Arithmetic_Logic_Unit.scala 171:58:@556.4]
  wire  _T_508; // @[Arithmetic_Logic_Unit.scala 171:58:@557.4]
  wire  _T_509; // @[Arithmetic_Logic_Unit.scala 171:58:@558.4]
  wire  _T_510; // @[Arithmetic_Logic_Unit.scala 171:58:@559.4]
  wire  _T_511; // @[Arithmetic_Logic_Unit.scala 171:58:@560.4]
  wire  _T_512; // @[Arithmetic_Logic_Unit.scala 171:58:@561.4]
  wire  _T_513; // @[Arithmetic_Logic_Unit.scala 171:58:@562.4]
  wire  _T_516; // @[Arithmetic_Logic_Unit.scala 171:55:@564.4]
  wire  _T_517; // @[Arithmetic_Logic_Unit.scala 171:55:@565.4]
  wire  _T_518; // @[Arithmetic_Logic_Unit.scala 171:55:@566.4]
  wire  _T_519; // @[Arithmetic_Logic_Unit.scala 171:55:@567.4]
  wire  _T_520; // @[Arithmetic_Logic_Unit.scala 171:55:@568.4]
  wire  _T_521; // @[Arithmetic_Logic_Unit.scala 171:55:@569.4]
  wire  _T_522; // @[Arithmetic_Logic_Unit.scala 171:55:@570.4]
  wire  _T_523; // @[Arithmetic_Logic_Unit.scala 171:55:@571.4]
  wire  _T_524; // @[Arithmetic_Logic_Unit.scala 171:55:@572.4]
  wire  _T_525; // @[Arithmetic_Logic_Unit.scala 171:55:@573.4]
  wire  _T_526; // @[Arithmetic_Logic_Unit.scala 171:55:@574.4]
  wire  _T_527; // @[Arithmetic_Logic_Unit.scala 171:55:@575.4]
  wire  _T_528; // @[Arithmetic_Logic_Unit.scala 171:55:@576.4]
  wire  _T_529; // @[Arithmetic_Logic_Unit.scala 171:55:@577.4]
  wire  _T_530; // @[Arithmetic_Logic_Unit.scala 171:55:@578.4]
  wire  _T_531; // @[Arithmetic_Logic_Unit.scala 171:55:@579.4]
  wire  _T_532; // @[Arithmetic_Logic_Unit.scala 171:55:@580.4]
  wire  _T_533; // @[Arithmetic_Logic_Unit.scala 171:55:@581.4]
  wire  _T_534; // @[Arithmetic_Logic_Unit.scala 171:55:@582.4]
  wire  _T_535; // @[Arithmetic_Logic_Unit.scala 171:55:@583.4]
  wire  _T_536; // @[Arithmetic_Logic_Unit.scala 171:55:@584.4]
  wire  _T_537; // @[Arithmetic_Logic_Unit.scala 171:55:@585.4]
  wire  _T_538; // @[Arithmetic_Logic_Unit.scala 171:55:@586.4]
  wire  _T_539; // @[Arithmetic_Logic_Unit.scala 171:55:@587.4]
  wire  _T_540; // @[Arithmetic_Logic_Unit.scala 171:55:@588.4]
  wire  _T_541; // @[Arithmetic_Logic_Unit.scala 171:55:@589.4]
  wire  _T_542; // @[Arithmetic_Logic_Unit.scala 171:55:@590.4]
  wire  _T_543; // @[Arithmetic_Logic_Unit.scala 171:55:@591.4]
  wire  _T_544; // @[Arithmetic_Logic_Unit.scala 171:55:@592.4]
  wire  _T_545; // @[Arithmetic_Logic_Unit.scala 171:55:@593.4]
  wire [31:0] result_unsigned; // @[Arithmetic_Logic_Unit.scala 65:29:@113.4 Arithmetic_Logic_Unit.scala 66:40:@115.4 Arithmetic_Logic_Unit.scala 78:19:@126.4 Arithmetic_Logic_Unit.scala 95:82:@132.6 Arithmetic_Logic_Unit.scala 96:82:@136.6 Arithmetic_Logic_Unit.scala 97:82:@142.6 Arithmetic_Logic_Unit.scala 98:82:@149.6 Arithmetic_Logic_Unit.scala 99:82:@155.6 Arithmetic_Logic_Unit.scala 100:82:@160.6 Arithmetic_Logic_Unit.scala 101:80:@165.6 Arithmetic_Logic_Unit.scala 102:80:@170.6 Arithmetic_Logic_Unit.scala 103:82:@175.6 Arithmetic_Logic_Unit.scala 104:83:@180.6 Arithmetic_Logic_Unit.scala 105:82:@185.6 Arithmetic_Logic_Unit.scala 106:82:@190.6 Arithmetic_Logic_Unit.scala 107:84:@195.6 Arithmetic_Logic_Unit.scala 108:86:@201.6 Arithmetic_Logic_Unit.scala 109:82:@206.6 Arithmetic_Logic_Unit.scala 110:84:@212.6 Arithmetic_Logic_Unit.scala 111:84:@217.6 Arithmetic_Logic_Unit.scala 112:86:@223.6 Arithmetic_Logic_Unit.scala 113:84:@228.6 Arithmetic_Logic_Unit.scala 114:86:@234.6 Arithmetic_Logic_Unit.scala 115:82:@239.6 Arithmetic_Logic_Unit.scala 116:84:@245.6 Arithmetic_Logic_Unit.scala 117:84:@252.6 Arithmetic_Logic_Unit.scala 118:86:@260.6 Arithmetic_Logic_Unit.scala 119:80:@266.6 Arithmetic_Logic_Unit.scala 122:25:@274.8 Arithmetic_Logic_Unit.scala 124:25:@281.8 Arithmetic_Logic_Unit.scala 127:80:@290.6 Arithmetic_Logic_Unit.scala 128:80:@297.6 Arithmetic_Logic_Unit.scala 131:25:@303.8 Arithmetic_Logic_Unit.scala 133:25:@418.8 Arithmetic_Logic_Unit.scala 138:25:@425.8 Arithmetic_Logic_Unit.scala 140:25:@491.8 Arithmetic_Logic_Unit.scala 144:23:@496.6]
  wire  _T_636; // @[Arithmetic_Logic_Unit.scala 181:9:@666.4]
  assign logical_operand0_unsigned = io_0 != 32'h0; // @[Arithmetic_Logic_Unit.scala 91:58:@127.4]
  assign logical_operand1_unsigned = io_1 != 32'h0; // @[Arithmetic_Logic_Unit.scala 92:58:@128.4]
  assign logical_operand2_unsigned = io_3 != 32'h0; // @[Arithmetic_Logic_Unit.scala 93:58:@129.4]
  assign _T_43 = io_4 == 5'h1; // @[Arithmetic_Logic_Unit.scala 96:49:@134.4]
  assign _GEN_1 = _T_43 ? io_0 : 32'h0; // @[Arithmetic_Logic_Unit.scala 96:65:@135.4]
  assign _T_45 = io_4 == 5'h2; // @[Arithmetic_Logic_Unit.scala 97:49:@138.4]
  assign _T_46 = io_0 + io_1; // @[Arithmetic_Logic_Unit.scala 97:103:@140.6]
  assign _T_47 = io_0 + io_1; // @[Arithmetic_Logic_Unit.scala 97:103:@141.6]
  assign _GEN_2 = _T_45 ? _T_47 : _GEN_1; // @[Arithmetic_Logic_Unit.scala 97:65:@139.4]
  assign _T_49 = io_4 == 5'h3; // @[Arithmetic_Logic_Unit.scala 98:49:@144.4]
  assign _T_50 = io_0 - io_1; // @[Arithmetic_Logic_Unit.scala 98:103:@146.6]
  assign _T_51 = $unsigned(_T_50); // @[Arithmetic_Logic_Unit.scala 98:103:@147.6]
  assign _T_52 = _T_51[31:0]; // @[Arithmetic_Logic_Unit.scala 98:103:@148.6]
  assign _GEN_3 = _T_49 ? _T_52 : _GEN_2; // @[Arithmetic_Logic_Unit.scala 98:65:@145.4]
  assign _T_54 = io_4 == 5'h4; // @[Arithmetic_Logic_Unit.scala 99:49:@151.4]
  assign _T_55 = io_1[18:0]; // @[Arithmetic_Logic_Unit.scala 99:123:@153.6]
  assign _GEN_37 = {{524287'd0}, io_0}; // @[Arithmetic_Logic_Unit.scala 99:103:@154.6]
  assign _T_56 = _GEN_37 << _T_55; // @[Arithmetic_Logic_Unit.scala 99:103:@154.6]
  assign _GEN_4 = _T_54 ? _T_56 : {{524287'd0}, _GEN_3}; // @[Arithmetic_Logic_Unit.scala 99:65:@152.4]
  assign _T_58 = io_4 == 5'h6; // @[Arithmetic_Logic_Unit.scala 100:49:@157.4]
  assign _T_59 = io_0 >> io_1; // @[Arithmetic_Logic_Unit.scala 100:103:@159.6]
  assign _GEN_5 = _T_58 ? {{524287'd0}, _T_59} : _GEN_4; // @[Arithmetic_Logic_Unit.scala 100:65:@158.4]
  assign _T_61 = io_4 == 5'h7; // @[Arithmetic_Logic_Unit.scala 101:48:@162.4]
  assign _T_62 = io_0 == io_1; // @[Arithmetic_Logic_Unit.scala 101:101:@164.6]
  assign _GEN_6 = _T_61 ? {{524318'd0}, _T_62} : _GEN_5; // @[Arithmetic_Logic_Unit.scala 101:63:@163.4]
  assign _T_64 = io_4 == 5'h8; // @[Arithmetic_Logic_Unit.scala 102:48:@167.4]
  assign _T_65 = io_0 != io_1; // @[Arithmetic_Logic_Unit.scala 102:101:@169.6]
  assign _GEN_7 = _T_64 ? {{524318'd0}, _T_65} : _GEN_6; // @[Arithmetic_Logic_Unit.scala 102:63:@168.4]
  assign _T_67 = io_4 == 5'ha; // @[Arithmetic_Logic_Unit.scala 103:49:@172.4]
  assign _T_68 = io_0 > io_1; // @[Arithmetic_Logic_Unit.scala 103:103:@174.6]
  assign _GEN_8 = _T_67 ? {{524318'd0}, _T_68} : _GEN_7; // @[Arithmetic_Logic_Unit.scala 103:65:@173.4]
  assign _T_70 = io_4 == 5'hc; // @[Arithmetic_Logic_Unit.scala 104:49:@177.4]
  assign _T_71 = io_0 < io_1; // @[Arithmetic_Logic_Unit.scala 104:104:@179.6]
  assign _GEN_9 = _T_70 ? {{524318'd0}, _T_71} : _GEN_8; // @[Arithmetic_Logic_Unit.scala 104:66:@178.4]
  assign _T_73 = io_4 == 5'he; // @[Arithmetic_Logic_Unit.scala 105:49:@182.4]
  assign _T_74 = io_0 >= io_1; // @[Arithmetic_Logic_Unit.scala 105:103:@184.6]
  assign _GEN_10 = _T_73 ? {{524318'd0}, _T_74} : _GEN_9; // @[Arithmetic_Logic_Unit.scala 105:65:@183.4]
  assign _T_76 = io_4 == 5'h10; // @[Arithmetic_Logic_Unit.scala 106:49:@187.4]
  assign _T_77 = io_0 <= io_1; // @[Arithmetic_Logic_Unit.scala 106:103:@189.6]
  assign _GEN_11 = _T_76 ? {{524318'd0}, _T_77} : _GEN_10; // @[Arithmetic_Logic_Unit.scala 106:65:@188.4]
  assign _T_79 = io_4 == 5'h11; // @[Arithmetic_Logic_Unit.scala 107:50:@192.4]
  assign _T_80 = io_0 & io_1; // @[Arithmetic_Logic_Unit.scala 107:105:@194.6]
  assign _GEN_12 = _T_79 ? {{524287'd0}, _T_80} : _GEN_11; // @[Arithmetic_Logic_Unit.scala 107:67:@193.4]
  assign _T_82 = io_4 == 5'h12; // @[Arithmetic_Logic_Unit.scala 108:51:@197.4]
  assign _T_84 = ~ _T_80; // @[Arithmetic_Logic_Unit.scala 108:89:@200.6]
  assign _GEN_13 = _T_82 ? {{524287'd0}, _T_84} : _GEN_12; // @[Arithmetic_Logic_Unit.scala 108:69:@198.4]
  assign _T_86 = io_4 == 5'h13; // @[Arithmetic_Logic_Unit.scala 109:49:@203.4]
  assign _T_87 = io_0 | io_1; // @[Arithmetic_Logic_Unit.scala 109:103:@205.6]
  assign _GEN_14 = _T_86 ? {{524287'd0}, _T_87} : _GEN_13; // @[Arithmetic_Logic_Unit.scala 109:65:@204.4]
  assign _T_89 = io_4 == 5'h14; // @[Arithmetic_Logic_Unit.scala 110:50:@208.4]
  assign _T_91 = ~ _T_87; // @[Arithmetic_Logic_Unit.scala 110:87:@211.6]
  assign _GEN_15 = _T_89 ? {{524287'd0}, _T_91} : _GEN_14; // @[Arithmetic_Logic_Unit.scala 110:67:@209.4]
  assign _T_93 = io_4 == 5'h15; // @[Arithmetic_Logic_Unit.scala 111:50:@214.4]
  assign _T_94 = io_0 ^ io_1; // @[Arithmetic_Logic_Unit.scala 111:105:@216.6]
  assign _GEN_16 = _T_93 ? {{524287'd0}, _T_94} : _GEN_15; // @[Arithmetic_Logic_Unit.scala 111:67:@215.4]
  assign _T_96 = io_4 == 5'h16; // @[Arithmetic_Logic_Unit.scala 112:51:@219.4]
  assign _T_98 = ~ _T_94; // @[Arithmetic_Logic_Unit.scala 112:89:@222.6]
  assign _GEN_17 = _T_96 ? {{524287'd0}, _T_98} : _GEN_16; // @[Arithmetic_Logic_Unit.scala 112:69:@220.4]
  assign _T_100 = io_4 == 5'h17; // @[Arithmetic_Logic_Unit.scala 113:50:@225.4]
  assign _T_101 = logical_operand0_unsigned & logical_operand1_unsigned; // @[Arithmetic_Logic_Unit.scala 113:113:@227.6]
  assign _GEN_18 = _T_100 ? {{524318'd0}, _T_101} : _GEN_17; // @[Arithmetic_Logic_Unit.scala 113:67:@226.4]
  assign _T_103 = io_4 == 5'h18; // @[Arithmetic_Logic_Unit.scala 114:51:@230.4]
  assign _T_106 = _T_101 == 1'h0; // @[Arithmetic_Logic_Unit.scala 114:89:@233.6]
  assign _GEN_19 = _T_103 ? {{524318'd0}, _T_106} : _GEN_18; // @[Arithmetic_Logic_Unit.scala 114:69:@231.4]
  assign _T_108 = io_4 == 5'h19; // @[Arithmetic_Logic_Unit.scala 115:49:@236.4]
  assign _T_109 = logical_operand0_unsigned | logical_operand1_unsigned; // @[Arithmetic_Logic_Unit.scala 115:111:@238.6]
  assign _GEN_20 = _T_108 ? {{524318'd0}, _T_109} : _GEN_19; // @[Arithmetic_Logic_Unit.scala 115:65:@237.4]
  assign _T_111 = io_4 == 5'h1a; // @[Arithmetic_Logic_Unit.scala 116:50:@241.4]
  assign _T_114 = _T_109 == 1'h0; // @[Arithmetic_Logic_Unit.scala 116:87:@244.6]
  assign _GEN_21 = _T_111 ? {{524318'd0}, _T_114} : _GEN_20; // @[Arithmetic_Logic_Unit.scala 116:67:@242.4]
  assign _T_116 = io_4 == 5'h1b; // @[Arithmetic_Logic_Unit.scala 117:50:@247.4]
  assign _T_118 = logical_operand0_unsigned == 1'h0; // @[Arithmetic_Logic_Unit.scala 117:87:@249.6]
  assign _T_120 = logical_operand1_unsigned == 1'h0; // @[Arithmetic_Logic_Unit.scala 117:116:@250.6]
  assign _T_121 = _T_118 ^ _T_120; // @[Arithmetic_Logic_Unit.scala 117:114:@251.6]
  assign _GEN_22 = _T_116 ? {{524318'd0}, _T_121} : _GEN_21; // @[Arithmetic_Logic_Unit.scala 117:67:@248.4]
  assign _T_123 = io_4 == 5'h1c; // @[Arithmetic_Logic_Unit.scala 118:51:@254.4]
  assign _T_130 = _T_121 == 1'h0; // @[Arithmetic_Logic_Unit.scala 118:89:@259.6]
  assign _GEN_23 = _T_123 ? {{524318'd0}, _T_130} : _GEN_22; // @[Arithmetic_Logic_Unit.scala 118:69:@255.4]
  assign _GEN_38 = {{1'd0}, io_4}; // @[Arithmetic_Logic_Unit.scala 119:48:@262.4]
  assign _T_132 = _GEN_38 == 6'h21; // @[Arithmetic_Logic_Unit.scala 119:48:@262.4]
  assign _T_134 = _T_59[0]; // @[Arithmetic_Logic_Unit.scala 119:100:@265.6]
  assign _GEN_24 = _T_132 ? {{524318'd0}, _T_134} : _GEN_23; // @[Arithmetic_Logic_Unit.scala 119:63:@263.4]
  assign _T_136 = _GEN_38 == 6'h22; // @[Arithmetic_Logic_Unit.scala 120:48:@268.4]
  assign _T_139 = 524288'h1 << _T_55; // @[Arithmetic_Logic_Unit.scala 122:53:@272.8]
  assign _GEN_40 = {{524256'd0}, io_0}; // @[Arithmetic_Logic_Unit.scala 122:46:@273.8]
  assign _T_140 = _GEN_40 | _T_139; // @[Arithmetic_Logic_Unit.scala 122:46:@273.8]
  assign _T_144 = ~ _T_139; // @[Arithmetic_Logic_Unit.scala 124:49:@279.8]
  assign _T_145 = _GEN_40 & _T_144; // @[Arithmetic_Logic_Unit.scala 124:46:@280.8]
  assign _GEN_25 = logical_operand2_unsigned ? _T_140 : _T_145; // @[Arithmetic_Logic_Unit.scala 121:38:@270.6]
  assign _GEN_26 = _T_136 ? {{31'd0}, _GEN_25} : _GEN_24; // @[Arithmetic_Logic_Unit.scala 120:63:@269.4]
  assign _T_147 = _GEN_38 == 6'h23; // @[Arithmetic_Logic_Unit.scala 127:48:@284.4]
  assign _GEN_27 = _T_147 ? {{31'd0}, _T_145} : _GEN_26; // @[Arithmetic_Logic_Unit.scala 127:63:@285.4]
  assign _T_154 = _GEN_38 == 6'h24; // @[Arithmetic_Logic_Unit.scala 128:48:@292.4]
  assign _GEN_28 = _T_154 ? {{31'd0}, _T_140} : _GEN_27; // @[Arithmetic_Logic_Unit.scala 128:63:@293.4]
  assign _T_160 = _GEN_38 == 6'h25; // @[Arithmetic_Logic_Unit.scala 129:49:@299.4]
  assign _T_162 = io_0 == 32'h0; // @[Arithmetic_Logic_Unit.scala 130:30:@301.6]
  assign _T_168 = io_0[31:16]; // @[Bitwise.scala 103:21:@308.8]
  assign _T_169 = {{16'd0}, _T_168}; // @[Bitwise.scala 103:31:@309.8]
  assign _T_170 = io_0[15:0]; // @[Bitwise.scala 103:46:@310.8]
  assign _GEN_47 = {{16'd0}, _T_170}; // @[Bitwise.scala 103:65:@311.8]
  assign _T_171 = _GEN_47 << 16; // @[Bitwise.scala 103:65:@311.8]
  assign _T_173 = _T_171 & 32'hffff0000; // @[Bitwise.scala 103:75:@313.8]
  assign _T_174 = _T_169 | _T_173; // @[Bitwise.scala 103:39:@314.8]
  assign _T_178 = _T_174[31:8]; // @[Bitwise.scala 103:21:@318.8]
  assign _GEN_48 = {{8'd0}, _T_178}; // @[Bitwise.scala 103:31:@319.8]
  assign _T_179 = _GEN_48 & 32'hff00ff; // @[Bitwise.scala 103:31:@319.8]
  assign _T_180 = _T_174[23:0]; // @[Bitwise.scala 103:46:@320.8]
  assign _GEN_49 = {{8'd0}, _T_180}; // @[Bitwise.scala 103:65:@321.8]
  assign _T_181 = _GEN_49 << 8; // @[Bitwise.scala 103:65:@321.8]
  assign _T_183 = _T_181 & 32'hff00ff00; // @[Bitwise.scala 103:75:@323.8]
  assign _T_184 = _T_179 | _T_183; // @[Bitwise.scala 103:39:@324.8]
  assign _T_188 = _T_184[31:4]; // @[Bitwise.scala 103:21:@328.8]
  assign _GEN_50 = {{4'd0}, _T_188}; // @[Bitwise.scala 103:31:@329.8]
  assign _T_189 = _GEN_50 & 32'hf0f0f0f; // @[Bitwise.scala 103:31:@329.8]
  assign _T_190 = _T_184[27:0]; // @[Bitwise.scala 103:46:@330.8]
  assign _GEN_51 = {{4'd0}, _T_190}; // @[Bitwise.scala 103:65:@331.8]
  assign _T_191 = _GEN_51 << 4; // @[Bitwise.scala 103:65:@331.8]
  assign _T_193 = _T_191 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75:@333.8]
  assign _T_194 = _T_189 | _T_193; // @[Bitwise.scala 103:39:@334.8]
  assign _T_198 = _T_194[31:2]; // @[Bitwise.scala 103:21:@338.8]
  assign _GEN_52 = {{2'd0}, _T_198}; // @[Bitwise.scala 103:31:@339.8]
  assign _T_199 = _GEN_52 & 32'h33333333; // @[Bitwise.scala 103:31:@339.8]
  assign _T_200 = _T_194[29:0]; // @[Bitwise.scala 103:46:@340.8]
  assign _GEN_53 = {{2'd0}, _T_200}; // @[Bitwise.scala 103:65:@341.8]
  assign _T_201 = _GEN_53 << 2; // @[Bitwise.scala 103:65:@341.8]
  assign _T_203 = _T_201 & 32'hcccccccc; // @[Bitwise.scala 103:75:@343.8]
  assign _T_204 = _T_199 | _T_203; // @[Bitwise.scala 103:39:@344.8]
  assign _T_208 = _T_204[31:1]; // @[Bitwise.scala 103:21:@348.8]
  assign _GEN_54 = {{1'd0}, _T_208}; // @[Bitwise.scala 103:31:@349.8]
  assign _T_209 = _GEN_54 & 32'h55555555; // @[Bitwise.scala 103:31:@349.8]
  assign _T_210 = _T_204[30:0]; // @[Bitwise.scala 103:46:@350.8]
  assign _GEN_55 = {{1'd0}, _T_210}; // @[Bitwise.scala 103:65:@351.8]
  assign _T_211 = _GEN_55 << 1; // @[Bitwise.scala 103:65:@351.8]
  assign _T_213 = _T_211 & 32'haaaaaaaa; // @[Bitwise.scala 103:75:@353.8]
  assign _T_214 = _T_209 | _T_213; // @[Bitwise.scala 103:39:@354.8]
  assign _T_215 = _T_214[0]; // @[OneHot.scala 39:40:@355.8]
  assign _T_216 = _T_214[1]; // @[OneHot.scala 39:40:@356.8]
  assign _T_217 = _T_214[2]; // @[OneHot.scala 39:40:@357.8]
  assign _T_218 = _T_214[3]; // @[OneHot.scala 39:40:@358.8]
  assign _T_219 = _T_214[4]; // @[OneHot.scala 39:40:@359.8]
  assign _T_220 = _T_214[5]; // @[OneHot.scala 39:40:@360.8]
  assign _T_221 = _T_214[6]; // @[OneHot.scala 39:40:@361.8]
  assign _T_222 = _T_214[7]; // @[OneHot.scala 39:40:@362.8]
  assign _T_223 = _T_214[8]; // @[OneHot.scala 39:40:@363.8]
  assign _T_224 = _T_214[9]; // @[OneHot.scala 39:40:@364.8]
  assign _T_225 = _T_214[10]; // @[OneHot.scala 39:40:@365.8]
  assign _T_226 = _T_214[11]; // @[OneHot.scala 39:40:@366.8]
  assign _T_227 = _T_214[12]; // @[OneHot.scala 39:40:@367.8]
  assign _T_228 = _T_214[13]; // @[OneHot.scala 39:40:@368.8]
  assign _T_229 = _T_214[14]; // @[OneHot.scala 39:40:@369.8]
  assign _T_230 = _T_214[15]; // @[OneHot.scala 39:40:@370.8]
  assign _T_231 = _T_214[16]; // @[OneHot.scala 39:40:@371.8]
  assign _T_232 = _T_214[17]; // @[OneHot.scala 39:40:@372.8]
  assign _T_233 = _T_214[18]; // @[OneHot.scala 39:40:@373.8]
  assign _T_234 = _T_214[19]; // @[OneHot.scala 39:40:@374.8]
  assign _T_235 = _T_214[20]; // @[OneHot.scala 39:40:@375.8]
  assign _T_236 = _T_214[21]; // @[OneHot.scala 39:40:@376.8]
  assign _T_237 = _T_214[22]; // @[OneHot.scala 39:40:@377.8]
  assign _T_238 = _T_214[23]; // @[OneHot.scala 39:40:@378.8]
  assign _T_239 = _T_214[24]; // @[OneHot.scala 39:40:@379.8]
  assign _T_240 = _T_214[25]; // @[OneHot.scala 39:40:@380.8]
  assign _T_241 = _T_214[26]; // @[OneHot.scala 39:40:@381.8]
  assign _T_242 = _T_214[27]; // @[OneHot.scala 39:40:@382.8]
  assign _T_243 = _T_214[28]; // @[OneHot.scala 39:40:@383.8]
  assign _T_244 = _T_214[29]; // @[OneHot.scala 39:40:@384.8]
  assign _T_245 = _T_214[30]; // @[OneHot.scala 39:40:@385.8]
  assign _T_279 = _T_245 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@387.8]
  assign _T_280 = _T_244 ? 5'h1d : _T_279; // @[Mux.scala 31:69:@388.8]
  assign _T_281 = _T_243 ? 5'h1c : _T_280; // @[Mux.scala 31:69:@389.8]
  assign _T_282 = _T_242 ? 5'h1b : _T_281; // @[Mux.scala 31:69:@390.8]
  assign _T_283 = _T_241 ? 5'h1a : _T_282; // @[Mux.scala 31:69:@391.8]
  assign _T_284 = _T_240 ? 5'h19 : _T_283; // @[Mux.scala 31:69:@392.8]
  assign _T_285 = _T_239 ? 5'h18 : _T_284; // @[Mux.scala 31:69:@393.8]
  assign _T_286 = _T_238 ? 5'h17 : _T_285; // @[Mux.scala 31:69:@394.8]
  assign _T_287 = _T_237 ? 5'h16 : _T_286; // @[Mux.scala 31:69:@395.8]
  assign _T_288 = _T_236 ? 5'h15 : _T_287; // @[Mux.scala 31:69:@396.8]
  assign _T_289 = _T_235 ? 5'h14 : _T_288; // @[Mux.scala 31:69:@397.8]
  assign _T_290 = _T_234 ? 5'h13 : _T_289; // @[Mux.scala 31:69:@398.8]
  assign _T_291 = _T_233 ? 5'h12 : _T_290; // @[Mux.scala 31:69:@399.8]
  assign _T_292 = _T_232 ? 5'h11 : _T_291; // @[Mux.scala 31:69:@400.8]
  assign _T_293 = _T_231 ? 5'h10 : _T_292; // @[Mux.scala 31:69:@401.8]
  assign _T_294 = _T_230 ? 5'hf : _T_293; // @[Mux.scala 31:69:@402.8]
  assign _T_295 = _T_229 ? 5'he : _T_294; // @[Mux.scala 31:69:@403.8]
  assign _T_296 = _T_228 ? 5'hd : _T_295; // @[Mux.scala 31:69:@404.8]
  assign _T_297 = _T_227 ? 5'hc : _T_296; // @[Mux.scala 31:69:@405.8]
  assign _T_298 = _T_226 ? 5'hb : _T_297; // @[Mux.scala 31:69:@406.8]
  assign _T_299 = _T_225 ? 5'ha : _T_298; // @[Mux.scala 31:69:@407.8]
  assign _T_300 = _T_224 ? 5'h9 : _T_299; // @[Mux.scala 31:69:@408.8]
  assign _T_301 = _T_223 ? 5'h8 : _T_300; // @[Mux.scala 31:69:@409.8]
  assign _T_302 = _T_222 ? 5'h7 : _T_301; // @[Mux.scala 31:69:@410.8]
  assign _T_303 = _T_221 ? 5'h6 : _T_302; // @[Mux.scala 31:69:@411.8]
  assign _T_304 = _T_220 ? 5'h5 : _T_303; // @[Mux.scala 31:69:@412.8]
  assign _T_305 = _T_219 ? 5'h4 : _T_304; // @[Mux.scala 31:69:@413.8]
  assign _T_306 = _T_218 ? 5'h3 : _T_305; // @[Mux.scala 31:69:@414.8]
  assign _T_307 = _T_217 ? 5'h2 : _T_306; // @[Mux.scala 31:69:@415.8]
  assign _T_308 = _T_216 ? 5'h1 : _T_307; // @[Mux.scala 31:69:@416.8]
  assign _T_309 = _T_215 ? 5'h0 : _T_308; // @[Mux.scala 31:69:@417.8]
  assign _GEN_29 = _T_162 ? 6'h20 : {{1'd0}, _T_309}; // @[Arithmetic_Logic_Unit.scala 130:38:@302.6]
  assign _GEN_30 = _T_160 ? {{524313'd0}, _GEN_29} : _GEN_28; // @[Arithmetic_Logic_Unit.scala 129:65:@300.4]
  assign _T_311 = _GEN_38 == 6'h26; // @[Arithmetic_Logic_Unit.scala 136:49:@421.4]
  assign _T_315 = io_0[0]; // @[OneHot.scala 39:40:@428.8]
  assign _T_316 = io_0[1]; // @[OneHot.scala 39:40:@429.8]
  assign _T_317 = io_0[2]; // @[OneHot.scala 39:40:@430.8]
  assign _T_318 = io_0[3]; // @[OneHot.scala 39:40:@431.8]
  assign _T_319 = io_0[4]; // @[OneHot.scala 39:40:@432.8]
  assign _T_320 = io_0[5]; // @[OneHot.scala 39:40:@433.8]
  assign _T_321 = io_0[6]; // @[OneHot.scala 39:40:@434.8]
  assign _T_322 = io_0[7]; // @[OneHot.scala 39:40:@435.8]
  assign _T_323 = io_0[8]; // @[OneHot.scala 39:40:@436.8]
  assign _T_324 = io_0[9]; // @[OneHot.scala 39:40:@437.8]
  assign _T_325 = io_0[10]; // @[OneHot.scala 39:40:@438.8]
  assign _T_326 = io_0[11]; // @[OneHot.scala 39:40:@439.8]
  assign _T_327 = io_0[12]; // @[OneHot.scala 39:40:@440.8]
  assign _T_328 = io_0[13]; // @[OneHot.scala 39:40:@441.8]
  assign _T_329 = io_0[14]; // @[OneHot.scala 39:40:@442.8]
  assign _T_330 = io_0[15]; // @[OneHot.scala 39:40:@443.8]
  assign _T_331 = io_0[16]; // @[OneHot.scala 39:40:@444.8]
  assign _T_332 = io_0[17]; // @[OneHot.scala 39:40:@445.8]
  assign _T_333 = io_0[18]; // @[OneHot.scala 39:40:@446.8]
  assign _T_334 = io_0[19]; // @[OneHot.scala 39:40:@447.8]
  assign _T_335 = io_0[20]; // @[OneHot.scala 39:40:@448.8]
  assign _T_336 = io_0[21]; // @[OneHot.scala 39:40:@449.8]
  assign _T_337 = io_0[22]; // @[OneHot.scala 39:40:@450.8]
  assign _T_338 = io_0[23]; // @[OneHot.scala 39:40:@451.8]
  assign _T_339 = io_0[24]; // @[OneHot.scala 39:40:@452.8]
  assign _T_340 = io_0[25]; // @[OneHot.scala 39:40:@453.8]
  assign _T_341 = io_0[26]; // @[OneHot.scala 39:40:@454.8]
  assign _T_342 = io_0[27]; // @[OneHot.scala 39:40:@455.8]
  assign _T_343 = io_0[28]; // @[OneHot.scala 39:40:@456.8]
  assign _T_344 = io_0[29]; // @[OneHot.scala 39:40:@457.8]
  assign _T_345 = io_0[30]; // @[OneHot.scala 39:40:@458.8]
  assign _T_379 = _T_345 ? 5'h1e : 5'h1f; // @[Mux.scala 31:69:@460.8]
  assign _T_380 = _T_344 ? 5'h1d : _T_379; // @[Mux.scala 31:69:@461.8]
  assign _T_381 = _T_343 ? 5'h1c : _T_380; // @[Mux.scala 31:69:@462.8]
  assign _T_382 = _T_342 ? 5'h1b : _T_381; // @[Mux.scala 31:69:@463.8]
  assign _T_383 = _T_341 ? 5'h1a : _T_382; // @[Mux.scala 31:69:@464.8]
  assign _T_384 = _T_340 ? 5'h19 : _T_383; // @[Mux.scala 31:69:@465.8]
  assign _T_385 = _T_339 ? 5'h18 : _T_384; // @[Mux.scala 31:69:@466.8]
  assign _T_386 = _T_338 ? 5'h17 : _T_385; // @[Mux.scala 31:69:@467.8]
  assign _T_387 = _T_337 ? 5'h16 : _T_386; // @[Mux.scala 31:69:@468.8]
  assign _T_388 = _T_336 ? 5'h15 : _T_387; // @[Mux.scala 31:69:@469.8]
  assign _T_389 = _T_335 ? 5'h14 : _T_388; // @[Mux.scala 31:69:@470.8]
  assign _T_390 = _T_334 ? 5'h13 : _T_389; // @[Mux.scala 31:69:@471.8]
  assign _T_391 = _T_333 ? 5'h12 : _T_390; // @[Mux.scala 31:69:@472.8]
  assign _T_392 = _T_332 ? 5'h11 : _T_391; // @[Mux.scala 31:69:@473.8]
  assign _T_393 = _T_331 ? 5'h10 : _T_392; // @[Mux.scala 31:69:@474.8]
  assign _T_394 = _T_330 ? 5'hf : _T_393; // @[Mux.scala 31:69:@475.8]
  assign _T_395 = _T_329 ? 5'he : _T_394; // @[Mux.scala 31:69:@476.8]
  assign _T_396 = _T_328 ? 5'hd : _T_395; // @[Mux.scala 31:69:@477.8]
  assign _T_397 = _T_327 ? 5'hc : _T_396; // @[Mux.scala 31:69:@478.8]
  assign _T_398 = _T_326 ? 5'hb : _T_397; // @[Mux.scala 31:69:@479.8]
  assign _T_399 = _T_325 ? 5'ha : _T_398; // @[Mux.scala 31:69:@480.8]
  assign _T_400 = _T_324 ? 5'h9 : _T_399; // @[Mux.scala 31:69:@481.8]
  assign _T_401 = _T_323 ? 5'h8 : _T_400; // @[Mux.scala 31:69:@482.8]
  assign _T_402 = _T_322 ? 5'h7 : _T_401; // @[Mux.scala 31:69:@483.8]
  assign _T_403 = _T_321 ? 5'h6 : _T_402; // @[Mux.scala 31:69:@484.8]
  assign _T_404 = _T_320 ? 5'h5 : _T_403; // @[Mux.scala 31:69:@485.8]
  assign _T_405 = _T_319 ? 5'h4 : _T_404; // @[Mux.scala 31:69:@486.8]
  assign _T_406 = _T_318 ? 5'h3 : _T_405; // @[Mux.scala 31:69:@487.8]
  assign _T_407 = _T_317 ? 5'h2 : _T_406; // @[Mux.scala 31:69:@488.8]
  assign _T_408 = _T_316 ? 5'h1 : _T_407; // @[Mux.scala 31:69:@489.8]
  assign _T_409 = _T_315 ? 5'h0 : _T_408; // @[Mux.scala 31:69:@490.8]
  assign _GEN_31 = _T_162 ? 6'h20 : {{1'd0}, _T_409}; // @[Arithmetic_Logic_Unit.scala 137:39:@424.6]
  assign _GEN_32 = _T_311 ? {{524313'd0}, _GEN_31} : _GEN_30; // @[Arithmetic_Logic_Unit.scala 136:65:@422.4]
  assign _T_411 = _GEN_38 == 6'h27; // @[Arithmetic_Logic_Unit.scala 143:50:@494.4]
  assign _GEN_33 = _T_411 ? 524319'h0 : _GEN_32; // @[Arithmetic_Logic_Unit.scala 143:67:@495.4]
  assign _T_483 = 6'h0 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@532.4]
  assign _T_484 = 6'h1 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@533.4]
  assign _T_485 = 6'h2 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@534.4]
  assign _T_486 = 6'h3 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@535.4]
  assign _T_487 = 6'h4 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@536.4]
  assign _T_488 = 6'h6 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@537.4]
  assign _T_489 = 6'h7 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@538.4]
  assign _T_490 = 6'h8 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@539.4]
  assign _T_491 = 6'ha == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@540.4]
  assign _T_492 = 6'hc == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@541.4]
  assign _T_493 = 6'he == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@542.4]
  assign _T_494 = 6'h10 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@543.4]
  assign _T_495 = 6'h11 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@544.4]
  assign _T_496 = 6'h12 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@545.4]
  assign _T_497 = 6'h13 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@546.4]
  assign _T_498 = 6'h14 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@547.4]
  assign _T_499 = 6'h15 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@548.4]
  assign _T_500 = 6'h16 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@549.4]
  assign _T_501 = 6'h17 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@550.4]
  assign _T_502 = 6'h18 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@551.4]
  assign _T_503 = 6'h19 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@552.4]
  assign _T_504 = 6'h1a == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@553.4]
  assign _T_505 = 6'h1b == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@554.4]
  assign _T_506 = 6'h1c == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@555.4]
  assign _T_507 = 6'h21 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@556.4]
  assign _T_508 = 6'h22 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@557.4]
  assign _T_509 = 6'h23 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@558.4]
  assign _T_510 = 6'h24 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@559.4]
  assign _T_511 = 6'h25 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@560.4]
  assign _T_512 = 6'h26 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@561.4]
  assign _T_513 = 6'h27 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@562.4]
  assign _T_516 = _T_483 | _T_484; // @[Arithmetic_Logic_Unit.scala 171:55:@564.4]
  assign _T_517 = _T_516 | _T_485; // @[Arithmetic_Logic_Unit.scala 171:55:@565.4]
  assign _T_518 = _T_517 | _T_486; // @[Arithmetic_Logic_Unit.scala 171:55:@566.4]
  assign _T_519 = _T_518 | _T_487; // @[Arithmetic_Logic_Unit.scala 171:55:@567.4]
  assign _T_520 = _T_519 | _T_488; // @[Arithmetic_Logic_Unit.scala 171:55:@568.4]
  assign _T_521 = _T_520 | _T_489; // @[Arithmetic_Logic_Unit.scala 171:55:@569.4]
  assign _T_522 = _T_521 | _T_490; // @[Arithmetic_Logic_Unit.scala 171:55:@570.4]
  assign _T_523 = _T_522 | _T_491; // @[Arithmetic_Logic_Unit.scala 171:55:@571.4]
  assign _T_524 = _T_523 | _T_492; // @[Arithmetic_Logic_Unit.scala 171:55:@572.4]
  assign _T_525 = _T_524 | _T_493; // @[Arithmetic_Logic_Unit.scala 171:55:@573.4]
  assign _T_526 = _T_525 | _T_494; // @[Arithmetic_Logic_Unit.scala 171:55:@574.4]
  assign _T_527 = _T_526 | _T_495; // @[Arithmetic_Logic_Unit.scala 171:55:@575.4]
  assign _T_528 = _T_527 | _T_496; // @[Arithmetic_Logic_Unit.scala 171:55:@576.4]
  assign _T_529 = _T_528 | _T_497; // @[Arithmetic_Logic_Unit.scala 171:55:@577.4]
  assign _T_530 = _T_529 | _T_498; // @[Arithmetic_Logic_Unit.scala 171:55:@578.4]
  assign _T_531 = _T_530 | _T_499; // @[Arithmetic_Logic_Unit.scala 171:55:@579.4]
  assign _T_532 = _T_531 | _T_500; // @[Arithmetic_Logic_Unit.scala 171:55:@580.4]
  assign _T_533 = _T_532 | _T_501; // @[Arithmetic_Logic_Unit.scala 171:55:@581.4]
  assign _T_534 = _T_533 | _T_502; // @[Arithmetic_Logic_Unit.scala 171:55:@582.4]
  assign _T_535 = _T_534 | _T_503; // @[Arithmetic_Logic_Unit.scala 171:55:@583.4]
  assign _T_536 = _T_535 | _T_504; // @[Arithmetic_Logic_Unit.scala 171:55:@584.4]
  assign _T_537 = _T_536 | _T_505; // @[Arithmetic_Logic_Unit.scala 171:55:@585.4]
  assign _T_538 = _T_537 | _T_506; // @[Arithmetic_Logic_Unit.scala 171:55:@586.4]
  assign _T_539 = _T_538 | _T_507; // @[Arithmetic_Logic_Unit.scala 171:55:@587.4]
  assign _T_540 = _T_539 | _T_508; // @[Arithmetic_Logic_Unit.scala 171:55:@588.4]
  assign _T_541 = _T_540 | _T_509; // @[Arithmetic_Logic_Unit.scala 171:55:@589.4]
  assign _T_542 = _T_541 | _T_510; // @[Arithmetic_Logic_Unit.scala 171:55:@590.4]
  assign _T_543 = _T_542 | _T_511; // @[Arithmetic_Logic_Unit.scala 171:55:@591.4]
  assign _T_544 = _T_543 | _T_512; // @[Arithmetic_Logic_Unit.scala 171:55:@592.4]
  assign _T_545 = _T_544 | _T_513; // @[Arithmetic_Logic_Unit.scala 171:55:@593.4]
  assign result_unsigned = _GEN_33[31:0]; // @[Arithmetic_Logic_Unit.scala 65:29:@113.4 Arithmetic_Logic_Unit.scala 66:40:@115.4 Arithmetic_Logic_Unit.scala 78:19:@126.4 Arithmetic_Logic_Unit.scala 95:82:@132.6 Arithmetic_Logic_Unit.scala 96:82:@136.6 Arithmetic_Logic_Unit.scala 97:82:@142.6 Arithmetic_Logic_Unit.scala 98:82:@149.6 Arithmetic_Logic_Unit.scala 99:82:@155.6 Arithmetic_Logic_Unit.scala 100:82:@160.6 Arithmetic_Logic_Unit.scala 101:80:@165.6 Arithmetic_Logic_Unit.scala 102:80:@170.6 Arithmetic_Logic_Unit.scala 103:82:@175.6 Arithmetic_Logic_Unit.scala 104:83:@180.6 Arithmetic_Logic_Unit.scala 105:82:@185.6 Arithmetic_Logic_Unit.scala 106:82:@190.6 Arithmetic_Logic_Unit.scala 107:84:@195.6 Arithmetic_Logic_Unit.scala 108:86:@201.6 Arithmetic_Logic_Unit.scala 109:82:@206.6 Arithmetic_Logic_Unit.scala 110:84:@212.6 Arithmetic_Logic_Unit.scala 111:84:@217.6 Arithmetic_Logic_Unit.scala 112:86:@223.6 Arithmetic_Logic_Unit.scala 113:84:@228.6 Arithmetic_Logic_Unit.scala 114:86:@234.6 Arithmetic_Logic_Unit.scala 115:82:@239.6 Arithmetic_Logic_Unit.scala 116:84:@245.6 Arithmetic_Logic_Unit.scala 117:84:@252.6 Arithmetic_Logic_Unit.scala 118:86:@260.6 Arithmetic_Logic_Unit.scala 119:80:@266.6 Arithmetic_Logic_Unit.scala 122:25:@274.8 Arithmetic_Logic_Unit.scala 124:25:@281.8 Arithmetic_Logic_Unit.scala 127:80:@290.6 Arithmetic_Logic_Unit.scala 128:80:@297.6 Arithmetic_Logic_Unit.scala 131:25:@303.8 Arithmetic_Logic_Unit.scala 133:25:@418.8 Arithmetic_Logic_Unit.scala 138:25:@425.8 Arithmetic_Logic_Unit.scala 140:25:@491.8 Arithmetic_Logic_Unit.scala 144:23:@496.6]
  assign _T_636 = reset == 1'h0; // @[Arithmetic_Logic_Unit.scala 181:9:@666.4]
  assign io_2 = _T_545 ? result_unsigned : 32'h0; // @[Arithmetic_Logic_Unit.scala 172:22:@595.6 Arithmetic_Logic_Unit.scala 174:22:@616.8 Arithmetic_Logic_Unit.scala 176:22:@660.10 Arithmetic_Logic_Unit.scala 178:22:@663.10]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_636) begin
          $fwrite(32'h80000002,"opcode = %d\n",io_4); // @[Arithmetic_Logic_Unit.scala 181:9:@668.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_636) begin
          $fwrite(32'h80000002,"operand 0 = %d\n",io_0); // @[Arithmetic_Logic_Unit.scala 182:9:@673.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_636) begin
          $fwrite(32'h80000002,"operand 1 = %d\n",io_1); // @[Arithmetic_Logic_Unit.scala 183:9:@678.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_636) begin
          $fwrite(32'h80000002,"result = %d\n",io_2); // @[Arithmetic_Logic_Unit.scala 184:9:@683.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_636) begin
          $fwrite(32'h80000002,"-----------------------------------\n"); // @[Arithmetic_Logic_Unit.scala 185:9:@688.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Delay_Pipe_Hw_6( // @[:@1379.2]
  input         clock, // @[:@1380.4]
  input         reset, // @[:@1381.4]
  input  [2:0]  io_2, // @[:@1382.4]
  output [15:0] io_1, // @[:@1382.4]
  input  [15:0] io_0 // @[:@1382.4]
);
  reg [2:0] head; // @[Delay_Pipe.scala 45:21:@1384.4]
  reg [31:0] _RAND_0;
  reg [2:0] tail; // @[Delay_Pipe.scala 46:21:@1385.4]
  reg [31:0] _RAND_1;
  reg [2:0] delay; // @[Delay_Pipe.scala 47:23:@1386.4]
  reg [31:0] _RAND_2;
  reg [15:0] fifo_0; // @[Delay_Pipe.scala 50:21:@1394.4]
  reg [31:0] _RAND_3;
  reg [15:0] fifo_1; // @[Delay_Pipe.scala 50:21:@1394.4]
  reg [31:0] _RAND_4;
  reg [15:0] fifo_2; // @[Delay_Pipe.scala 50:21:@1394.4]
  reg [31:0] _RAND_5;
  reg [15:0] fifo_3; // @[Delay_Pipe.scala 50:21:@1394.4]
  reg [31:0] _RAND_6;
  reg [15:0] fifo_4; // @[Delay_Pipe.scala 50:21:@1394.4]
  reg [31:0] _RAND_7;
  reg [15:0] fifo_5; // @[Delay_Pipe.scala 50:21:@1394.4]
  reg [31:0] _RAND_8;
  wire [15:0] _GEN_1; // @[Delay_Pipe.scala 53:12:@1395.4]
  wire [15:0] _GEN_2; // @[Delay_Pipe.scala 53:12:@1395.4]
  wire [15:0] _GEN_3; // @[Delay_Pipe.scala 53:12:@1395.4]
  wire [15:0] _GEN_4; // @[Delay_Pipe.scala 53:12:@1395.4]
  wire [15:0] _GEN_6; // @[Delay_Pipe.scala 54:14:@1396.4]
  wire [15:0] _GEN_7; // @[Delay_Pipe.scala 54:14:@1396.4]
  wire [15:0] _GEN_8; // @[Delay_Pipe.scala 54:14:@1396.4]
  wire [15:0] _GEN_9; // @[Delay_Pipe.scala 54:14:@1396.4]
  wire [15:0] _GEN_10; // @[Delay_Pipe.scala 54:14:@1396.4]
  wire [15:0] _GEN_11; // @[Delay_Pipe.scala 54:14:@1396.4]
  wire [3:0] _T_83; // @[Delay_Pipe.scala 55:16:@1397.4]
  wire [2:0] _T_84; // @[Delay_Pipe.scala 55:16:@1398.4]
  wire [3:0] _T_86; // @[Delay_Pipe.scala 56:16:@1400.4]
  wire [2:0] _T_87; // @[Delay_Pipe.scala 56:16:@1401.4]
  wire  _T_88; // @[Delay_Pipe.scala 59:15:@1403.4]
  wire [15:0] _GEN_12; // @[Delay_Pipe.scala 59:32:@1404.4]
  wire [15:0] _GEN_13; // @[Delay_Pipe.scala 59:32:@1404.4]
  wire [15:0] _GEN_14; // @[Delay_Pipe.scala 59:32:@1404.4]
  wire [15:0] _GEN_15; // @[Delay_Pipe.scala 59:32:@1404.4]
  wire [15:0] _GEN_16; // @[Delay_Pipe.scala 59:32:@1404.4]
  wire [15:0] _GEN_17; // @[Delay_Pipe.scala 59:32:@1404.4]
  wire [2:0] _GEN_18; // @[Delay_Pipe.scala 59:32:@1404.4]
  wire [2:0] _GEN_19; // @[Delay_Pipe.scala 59:32:@1404.4]
  assign _GEN_1 = 3'h1 == head ? fifo_1 : fifo_0; // @[Delay_Pipe.scala 53:12:@1395.4]
  assign _GEN_2 = 3'h2 == head ? fifo_2 : _GEN_1; // @[Delay_Pipe.scala 53:12:@1395.4]
  assign _GEN_3 = 3'h3 == head ? fifo_3 : _GEN_2; // @[Delay_Pipe.scala 53:12:@1395.4]
  assign _GEN_4 = 3'h4 == head ? fifo_4 : _GEN_3; // @[Delay_Pipe.scala 53:12:@1395.4]
  assign _GEN_6 = 3'h0 == tail ? io_0 : fifo_0; // @[Delay_Pipe.scala 54:14:@1396.4]
  assign _GEN_7 = 3'h1 == tail ? io_0 : fifo_1; // @[Delay_Pipe.scala 54:14:@1396.4]
  assign _GEN_8 = 3'h2 == tail ? io_0 : fifo_2; // @[Delay_Pipe.scala 54:14:@1396.4]
  assign _GEN_9 = 3'h3 == tail ? io_0 : fifo_3; // @[Delay_Pipe.scala 54:14:@1396.4]
  assign _GEN_10 = 3'h4 == tail ? io_0 : fifo_4; // @[Delay_Pipe.scala 54:14:@1396.4]
  assign _GEN_11 = 3'h5 == tail ? io_0 : fifo_5; // @[Delay_Pipe.scala 54:14:@1396.4]
  assign _T_83 = head + 3'h1; // @[Delay_Pipe.scala 55:16:@1397.4]
  assign _T_84 = head + 3'h1; // @[Delay_Pipe.scala 55:16:@1398.4]
  assign _T_86 = tail + 3'h1; // @[Delay_Pipe.scala 56:16:@1400.4]
  assign _T_87 = tail + 3'h1; // @[Delay_Pipe.scala 56:16:@1401.4]
  assign _T_88 = delay != io_2; // @[Delay_Pipe.scala 59:15:@1403.4]
  assign _GEN_12 = _T_88 ? 16'h0 : _GEN_6; // @[Delay_Pipe.scala 59:32:@1404.4]
  assign _GEN_13 = _T_88 ? 16'h0 : _GEN_7; // @[Delay_Pipe.scala 59:32:@1404.4]
  assign _GEN_14 = _T_88 ? 16'h0 : _GEN_8; // @[Delay_Pipe.scala 59:32:@1404.4]
  assign _GEN_15 = _T_88 ? 16'h0 : _GEN_9; // @[Delay_Pipe.scala 59:32:@1404.4]
  assign _GEN_16 = _T_88 ? 16'h0 : _GEN_10; // @[Delay_Pipe.scala 59:32:@1404.4]
  assign _GEN_17 = _T_88 ? 16'h0 : _GEN_11; // @[Delay_Pipe.scala 59:32:@1404.4]
  assign _GEN_18 = _T_88 ? io_2 : _T_87; // @[Delay_Pipe.scala 59:32:@1404.4]
  assign _GEN_19 = _T_88 ? io_2 : delay; // @[Delay_Pipe.scala 59:32:@1404.4]
  assign io_1 = 3'h5 == head ? fifo_5 : _GEN_4; // @[Delay_Pipe.scala 53:12:@1395.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  delay = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  fifo_0 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  fifo_1 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  fifo_2 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fifo_3 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  fifo_4 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  fifo_5 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      head <= 3'h0;
    end else begin
      head <= _T_84;
    end
    if (reset) begin
      tail <= 3'h0;
    end else begin
      if (_T_88) begin
        tail <= io_2;
      end else begin
        tail <= _T_87;
      end
    end
    if (reset) begin
      delay <= 3'h0;
    end else begin
      if (_T_88) begin
        delay <= io_2;
      end
    end
    if (reset) begin
      fifo_0 <= 16'h0;
    end else begin
      if (_T_88) begin
        fifo_0 <= 16'h0;
      end else begin
        if (3'h0 == tail) begin
          fifo_0 <= io_0;
        end
      end
    end
    if (reset) begin
      fifo_1 <= 16'h0;
    end else begin
      if (_T_88) begin
        fifo_1 <= 16'h0;
      end else begin
        if (3'h1 == tail) begin
          fifo_1 <= io_0;
        end
      end
    end
    if (reset) begin
      fifo_2 <= 16'h0;
    end else begin
      if (_T_88) begin
        fifo_2 <= 16'h0;
      end else begin
        if (3'h2 == tail) begin
          fifo_2 <= io_0;
        end
      end
    end
    if (reset) begin
      fifo_3 <= 16'h0;
    end else begin
      if (_T_88) begin
        fifo_3 <= 16'h0;
      end else begin
        if (3'h3 == tail) begin
          fifo_3 <= io_0;
        end
      end
    end
    if (reset) begin
      fifo_4 <= 16'h0;
    end else begin
      if (_T_88) begin
        fifo_4 <= 16'h0;
      end else begin
        if (3'h4 == tail) begin
          fifo_4 <= io_0;
        end
      end
    end
    if (reset) begin
      fifo_5 <= 16'h0;
    end else begin
      if (_T_88) begin
        fifo_5 <= 16'h0;
      end else begin
        if (3'h5 == tail) begin
          fifo_5 <= io_0;
        end
      end
    end
  end
endmodule
module Delay_Pipe_Hw_7( // @[:@1415.2]
  input         clock, // @[:@1416.4]
  input         reset, // @[:@1417.4]
  input  [1:0]  io_2, // @[:@1418.4]
  output [15:0] io_1, // @[:@1418.4]
  input  [15:0] io_0 // @[:@1418.4]
);
  reg [1:0] head; // @[Delay_Pipe.scala 45:21:@1420.4]
  reg [31:0] _RAND_0;
  reg [1:0] tail; // @[Delay_Pipe.scala 46:21:@1421.4]
  reg [31:0] _RAND_1;
  reg [1:0] delay; // @[Delay_Pipe.scala 47:23:@1422.4]
  reg [31:0] _RAND_2;
  reg [15:0] fifo_0; // @[Delay_Pipe.scala 50:21:@1427.4]
  reg [31:0] _RAND_3;
  reg [15:0] fifo_1; // @[Delay_Pipe.scala 50:21:@1427.4]
  reg [31:0] _RAND_4;
  reg [15:0] fifo_2; // @[Delay_Pipe.scala 50:21:@1427.4]
  reg [31:0] _RAND_5;
  wire [15:0] _GEN_1; // @[Delay_Pipe.scala 53:12:@1428.4]
  wire [15:0] _GEN_3; // @[Delay_Pipe.scala 54:14:@1429.4]
  wire [15:0] _GEN_4; // @[Delay_Pipe.scala 54:14:@1429.4]
  wire [15:0] _GEN_5; // @[Delay_Pipe.scala 54:14:@1429.4]
  wire [2:0] _T_62; // @[Delay_Pipe.scala 55:16:@1430.4]
  wire [1:0] _T_63; // @[Delay_Pipe.scala 55:16:@1431.4]
  wire [2:0] _T_65; // @[Delay_Pipe.scala 56:16:@1433.4]
  wire [1:0] _T_66; // @[Delay_Pipe.scala 56:16:@1434.4]
  wire  _T_67; // @[Delay_Pipe.scala 59:15:@1436.4]
  wire [15:0] _GEN_6; // @[Delay_Pipe.scala 59:32:@1437.4]
  wire [15:0] _GEN_7; // @[Delay_Pipe.scala 59:32:@1437.4]
  wire [15:0] _GEN_8; // @[Delay_Pipe.scala 59:32:@1437.4]
  wire [1:0] _GEN_9; // @[Delay_Pipe.scala 59:32:@1437.4]
  wire [1:0] _GEN_10; // @[Delay_Pipe.scala 59:32:@1437.4]
  assign _GEN_1 = 2'h1 == head ? fifo_1 : fifo_0; // @[Delay_Pipe.scala 53:12:@1428.4]
  assign _GEN_3 = 2'h0 == tail ? io_0 : fifo_0; // @[Delay_Pipe.scala 54:14:@1429.4]
  assign _GEN_4 = 2'h1 == tail ? io_0 : fifo_1; // @[Delay_Pipe.scala 54:14:@1429.4]
  assign _GEN_5 = 2'h2 == tail ? io_0 : fifo_2; // @[Delay_Pipe.scala 54:14:@1429.4]
  assign _T_62 = head + 2'h1; // @[Delay_Pipe.scala 55:16:@1430.4]
  assign _T_63 = head + 2'h1; // @[Delay_Pipe.scala 55:16:@1431.4]
  assign _T_65 = tail + 2'h1; // @[Delay_Pipe.scala 56:16:@1433.4]
  assign _T_66 = tail + 2'h1; // @[Delay_Pipe.scala 56:16:@1434.4]
  assign _T_67 = delay != io_2; // @[Delay_Pipe.scala 59:15:@1436.4]
  assign _GEN_6 = _T_67 ? 16'h0 : _GEN_3; // @[Delay_Pipe.scala 59:32:@1437.4]
  assign _GEN_7 = _T_67 ? 16'h0 : _GEN_4; // @[Delay_Pipe.scala 59:32:@1437.4]
  assign _GEN_8 = _T_67 ? 16'h0 : _GEN_5; // @[Delay_Pipe.scala 59:32:@1437.4]
  assign _GEN_9 = _T_67 ? io_2 : _T_66; // @[Delay_Pipe.scala 59:32:@1437.4]
  assign _GEN_10 = _T_67 ? io_2 : delay; // @[Delay_Pipe.scala 59:32:@1437.4]
  assign io_1 = 2'h2 == head ? fifo_2 : _GEN_1; // @[Delay_Pipe.scala 53:12:@1428.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  delay = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  fifo_0 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  fifo_1 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  fifo_2 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      head <= 2'h0;
    end else begin
      head <= _T_63;
    end
    if (reset) begin
      tail <= 2'h0;
    end else begin
      if (_T_67) begin
        tail <= io_2;
      end else begin
        tail <= _T_66;
      end
    end
    if (reset) begin
      delay <= 2'h0;
    end else begin
      if (_T_67) begin
        delay <= io_2;
      end
    end
    if (reset) begin
      fifo_0 <= 16'h0;
    end else begin
      if (_T_67) begin
        fifo_0 <= 16'h0;
      end else begin
        if (2'h0 == tail) begin
          fifo_0 <= io_0;
        end
      end
    end
    if (reset) begin
      fifo_1 <= 16'h0;
    end else begin
      if (_T_67) begin
        fifo_1 <= 16'h0;
      end else begin
        if (2'h1 == tail) begin
          fifo_1 <= io_0;
        end
      end
    end
    if (reset) begin
      fifo_2 <= 16'h0;
    end else begin
      if (_T_67) begin
        fifo_2 <= 16'h0;
      end else begin
        if (2'h2 == tail) begin
          fifo_2 <= io_0;
        end
      end
    end
  end
endmodule
module Arithmetic_Logic_Unit_Hw_2( // @[:@1475.2]
  input         clock, // @[:@1476.4]
  input         reset, // @[:@1477.4]
  input  [4:0]  io_4, // @[:@1478.4]
  input  [15:0] io_3, // @[:@1478.4]
  output [15:0] io_2, // @[:@1478.4]
  input  [15:0] io_1, // @[:@1478.4]
  input  [15:0] io_0 // @[:@1478.4]
);
  wire  logical_operand0_unsigned; // @[Arithmetic_Logic_Unit.scala 91:58:@1503.4]
  wire  logical_operand1_unsigned; // @[Arithmetic_Logic_Unit.scala 92:58:@1504.4]
  wire  logical_operand2_unsigned; // @[Arithmetic_Logic_Unit.scala 93:58:@1505.4]
  wire  _T_43; // @[Arithmetic_Logic_Unit.scala 96:49:@1510.4]
  wire [15:0] _GEN_1; // @[Arithmetic_Logic_Unit.scala 96:65:@1511.4]
  wire  _T_45; // @[Arithmetic_Logic_Unit.scala 97:49:@1514.4]
  wire [16:0] _T_46; // @[Arithmetic_Logic_Unit.scala 97:103:@1516.6]
  wire [15:0] _T_47; // @[Arithmetic_Logic_Unit.scala 97:103:@1517.6]
  wire [15:0] _GEN_2; // @[Arithmetic_Logic_Unit.scala 97:65:@1515.4]
  wire  _T_49; // @[Arithmetic_Logic_Unit.scala 98:49:@1520.4]
  wire [16:0] _T_50; // @[Arithmetic_Logic_Unit.scala 98:103:@1522.6]
  wire [16:0] _T_51; // @[Arithmetic_Logic_Unit.scala 98:103:@1523.6]
  wire [15:0] _T_52; // @[Arithmetic_Logic_Unit.scala 98:103:@1524.6]
  wire [15:0] _GEN_3; // @[Arithmetic_Logic_Unit.scala 98:65:@1521.4]
  wire  _T_54; // @[Arithmetic_Logic_Unit.scala 99:49:@1527.4]
  wire [65550:0] _GEN_37; // @[Arithmetic_Logic_Unit.scala 99:103:@1530.6]
  wire [65550:0] _T_56; // @[Arithmetic_Logic_Unit.scala 99:103:@1530.6]
  wire [65550:0] _GEN_4; // @[Arithmetic_Logic_Unit.scala 99:65:@1528.4]
  wire  _T_58; // @[Arithmetic_Logic_Unit.scala 100:49:@1533.4]
  wire [15:0] _T_59; // @[Arithmetic_Logic_Unit.scala 100:103:@1535.6]
  wire [65550:0] _GEN_5; // @[Arithmetic_Logic_Unit.scala 100:65:@1534.4]
  wire  _T_61; // @[Arithmetic_Logic_Unit.scala 101:48:@1538.4]
  wire  _T_62; // @[Arithmetic_Logic_Unit.scala 101:101:@1540.6]
  wire [65550:0] _GEN_6; // @[Arithmetic_Logic_Unit.scala 101:63:@1539.4]
  wire  _T_64; // @[Arithmetic_Logic_Unit.scala 102:48:@1543.4]
  wire  _T_65; // @[Arithmetic_Logic_Unit.scala 102:101:@1545.6]
  wire [65550:0] _GEN_7; // @[Arithmetic_Logic_Unit.scala 102:63:@1544.4]
  wire  _T_67; // @[Arithmetic_Logic_Unit.scala 103:49:@1548.4]
  wire  _T_68; // @[Arithmetic_Logic_Unit.scala 103:103:@1550.6]
  wire [65550:0] _GEN_8; // @[Arithmetic_Logic_Unit.scala 103:65:@1549.4]
  wire  _T_70; // @[Arithmetic_Logic_Unit.scala 104:49:@1553.4]
  wire  _T_71; // @[Arithmetic_Logic_Unit.scala 104:104:@1555.6]
  wire [65550:0] _GEN_9; // @[Arithmetic_Logic_Unit.scala 104:66:@1554.4]
  wire  _T_73; // @[Arithmetic_Logic_Unit.scala 105:49:@1558.4]
  wire  _T_74; // @[Arithmetic_Logic_Unit.scala 105:103:@1560.6]
  wire [65550:0] _GEN_10; // @[Arithmetic_Logic_Unit.scala 105:65:@1559.4]
  wire  _T_76; // @[Arithmetic_Logic_Unit.scala 106:49:@1563.4]
  wire  _T_77; // @[Arithmetic_Logic_Unit.scala 106:103:@1565.6]
  wire [65550:0] _GEN_11; // @[Arithmetic_Logic_Unit.scala 106:65:@1564.4]
  wire  _T_79; // @[Arithmetic_Logic_Unit.scala 107:50:@1568.4]
  wire [15:0] _T_80; // @[Arithmetic_Logic_Unit.scala 107:105:@1570.6]
  wire [65550:0] _GEN_12; // @[Arithmetic_Logic_Unit.scala 107:67:@1569.4]
  wire  _T_82; // @[Arithmetic_Logic_Unit.scala 108:51:@1573.4]
  wire [15:0] _T_84; // @[Arithmetic_Logic_Unit.scala 108:89:@1576.6]
  wire [65550:0] _GEN_13; // @[Arithmetic_Logic_Unit.scala 108:69:@1574.4]
  wire  _T_86; // @[Arithmetic_Logic_Unit.scala 109:49:@1579.4]
  wire [15:0] _T_87; // @[Arithmetic_Logic_Unit.scala 109:103:@1581.6]
  wire [65550:0] _GEN_14; // @[Arithmetic_Logic_Unit.scala 109:65:@1580.4]
  wire  _T_89; // @[Arithmetic_Logic_Unit.scala 110:50:@1584.4]
  wire [15:0] _T_91; // @[Arithmetic_Logic_Unit.scala 110:87:@1587.6]
  wire [65550:0] _GEN_15; // @[Arithmetic_Logic_Unit.scala 110:67:@1585.4]
  wire  _T_93; // @[Arithmetic_Logic_Unit.scala 111:50:@1590.4]
  wire [15:0] _T_94; // @[Arithmetic_Logic_Unit.scala 111:105:@1592.6]
  wire [65550:0] _GEN_16; // @[Arithmetic_Logic_Unit.scala 111:67:@1591.4]
  wire  _T_96; // @[Arithmetic_Logic_Unit.scala 112:51:@1595.4]
  wire [15:0] _T_98; // @[Arithmetic_Logic_Unit.scala 112:89:@1598.6]
  wire [65550:0] _GEN_17; // @[Arithmetic_Logic_Unit.scala 112:69:@1596.4]
  wire  _T_100; // @[Arithmetic_Logic_Unit.scala 113:50:@1601.4]
  wire  _T_101; // @[Arithmetic_Logic_Unit.scala 113:113:@1603.6]
  wire [65550:0] _GEN_18; // @[Arithmetic_Logic_Unit.scala 113:67:@1602.4]
  wire  _T_103; // @[Arithmetic_Logic_Unit.scala 114:51:@1606.4]
  wire  _T_106; // @[Arithmetic_Logic_Unit.scala 114:89:@1609.6]
  wire [65550:0] _GEN_19; // @[Arithmetic_Logic_Unit.scala 114:69:@1607.4]
  wire  _T_108; // @[Arithmetic_Logic_Unit.scala 115:49:@1612.4]
  wire  _T_109; // @[Arithmetic_Logic_Unit.scala 115:111:@1614.6]
  wire [65550:0] _GEN_20; // @[Arithmetic_Logic_Unit.scala 115:65:@1613.4]
  wire  _T_111; // @[Arithmetic_Logic_Unit.scala 116:50:@1617.4]
  wire  _T_114; // @[Arithmetic_Logic_Unit.scala 116:87:@1620.6]
  wire [65550:0] _GEN_21; // @[Arithmetic_Logic_Unit.scala 116:67:@1618.4]
  wire  _T_116; // @[Arithmetic_Logic_Unit.scala 117:50:@1623.4]
  wire  _T_118; // @[Arithmetic_Logic_Unit.scala 117:87:@1625.6]
  wire  _T_120; // @[Arithmetic_Logic_Unit.scala 117:116:@1626.6]
  wire  _T_121; // @[Arithmetic_Logic_Unit.scala 117:114:@1627.6]
  wire [65550:0] _GEN_22; // @[Arithmetic_Logic_Unit.scala 117:67:@1624.4]
  wire  _T_123; // @[Arithmetic_Logic_Unit.scala 118:51:@1630.4]
  wire  _T_130; // @[Arithmetic_Logic_Unit.scala 118:89:@1635.6]
  wire [65550:0] _GEN_23; // @[Arithmetic_Logic_Unit.scala 118:69:@1631.4]
  wire [5:0] _GEN_38; // @[Arithmetic_Logic_Unit.scala 119:48:@1638.4]
  wire  _T_132; // @[Arithmetic_Logic_Unit.scala 119:48:@1638.4]
  wire  _T_134; // @[Arithmetic_Logic_Unit.scala 119:100:@1641.6]
  wire [65550:0] _GEN_24; // @[Arithmetic_Logic_Unit.scala 119:63:@1639.4]
  wire  _T_136; // @[Arithmetic_Logic_Unit.scala 120:48:@1644.4]
  wire [65535:0] _T_139; // @[Arithmetic_Logic_Unit.scala 122:53:@1648.8]
  wire [65535:0] _GEN_40; // @[Arithmetic_Logic_Unit.scala 122:46:@1649.8]
  wire [65535:0] _T_140; // @[Arithmetic_Logic_Unit.scala 122:46:@1649.8]
  wire [65535:0] _T_144; // @[Arithmetic_Logic_Unit.scala 124:49:@1655.8]
  wire [65535:0] _T_145; // @[Arithmetic_Logic_Unit.scala 124:46:@1656.8]
  wire [65535:0] _GEN_25; // @[Arithmetic_Logic_Unit.scala 121:38:@1646.6]
  wire [65550:0] _GEN_26; // @[Arithmetic_Logic_Unit.scala 120:63:@1645.4]
  wire  _T_147; // @[Arithmetic_Logic_Unit.scala 127:48:@1660.4]
  wire [65550:0] _GEN_27; // @[Arithmetic_Logic_Unit.scala 127:63:@1661.4]
  wire  _T_154; // @[Arithmetic_Logic_Unit.scala 128:48:@1668.4]
  wire [65550:0] _GEN_28; // @[Arithmetic_Logic_Unit.scala 128:63:@1669.4]
  wire  _T_160; // @[Arithmetic_Logic_Unit.scala 129:49:@1675.4]
  wire  _T_162; // @[Arithmetic_Logic_Unit.scala 130:30:@1677.6]
  wire [7:0] _T_168; // @[Bitwise.scala 103:21:@1684.8]
  wire [15:0] _T_169; // @[Bitwise.scala 103:31:@1685.8]
  wire [7:0] _T_170; // @[Bitwise.scala 103:46:@1686.8]
  wire [15:0] _GEN_47; // @[Bitwise.scala 103:65:@1687.8]
  wire [15:0] _T_171; // @[Bitwise.scala 103:65:@1687.8]
  wire [15:0] _T_173; // @[Bitwise.scala 103:75:@1689.8]
  wire [15:0] _T_174; // @[Bitwise.scala 103:39:@1690.8]
  wire [11:0] _T_178; // @[Bitwise.scala 103:21:@1694.8]
  wire [15:0] _GEN_48; // @[Bitwise.scala 103:31:@1695.8]
  wire [15:0] _T_179; // @[Bitwise.scala 103:31:@1695.8]
  wire [11:0] _T_180; // @[Bitwise.scala 103:46:@1696.8]
  wire [15:0] _GEN_49; // @[Bitwise.scala 103:65:@1697.8]
  wire [15:0] _T_181; // @[Bitwise.scala 103:65:@1697.8]
  wire [15:0] _T_183; // @[Bitwise.scala 103:75:@1699.8]
  wire [15:0] _T_184; // @[Bitwise.scala 103:39:@1700.8]
  wire [13:0] _T_188; // @[Bitwise.scala 103:21:@1704.8]
  wire [15:0] _GEN_50; // @[Bitwise.scala 103:31:@1705.8]
  wire [15:0] _T_189; // @[Bitwise.scala 103:31:@1705.8]
  wire [13:0] _T_190; // @[Bitwise.scala 103:46:@1706.8]
  wire [15:0] _GEN_51; // @[Bitwise.scala 103:65:@1707.8]
  wire [15:0] _T_191; // @[Bitwise.scala 103:65:@1707.8]
  wire [15:0] _T_193; // @[Bitwise.scala 103:75:@1709.8]
  wire [15:0] _T_194; // @[Bitwise.scala 103:39:@1710.8]
  wire [14:0] _T_198; // @[Bitwise.scala 103:21:@1714.8]
  wire [15:0] _GEN_52; // @[Bitwise.scala 103:31:@1715.8]
  wire [15:0] _T_199; // @[Bitwise.scala 103:31:@1715.8]
  wire [14:0] _T_200; // @[Bitwise.scala 103:46:@1716.8]
  wire [15:0] _GEN_53; // @[Bitwise.scala 103:65:@1717.8]
  wire [15:0] _T_201; // @[Bitwise.scala 103:65:@1717.8]
  wire [15:0] _T_203; // @[Bitwise.scala 103:75:@1719.8]
  wire [15:0] _T_204; // @[Bitwise.scala 103:39:@1720.8]
  wire  _T_205; // @[OneHot.scala 39:40:@1721.8]
  wire  _T_206; // @[OneHot.scala 39:40:@1722.8]
  wire  _T_207; // @[OneHot.scala 39:40:@1723.8]
  wire  _T_208; // @[OneHot.scala 39:40:@1724.8]
  wire  _T_209; // @[OneHot.scala 39:40:@1725.8]
  wire  _T_210; // @[OneHot.scala 39:40:@1726.8]
  wire  _T_211; // @[OneHot.scala 39:40:@1727.8]
  wire  _T_212; // @[OneHot.scala 39:40:@1728.8]
  wire  _T_213; // @[OneHot.scala 39:40:@1729.8]
  wire  _T_214; // @[OneHot.scala 39:40:@1730.8]
  wire  _T_215; // @[OneHot.scala 39:40:@1731.8]
  wire  _T_216; // @[OneHot.scala 39:40:@1732.8]
  wire  _T_217; // @[OneHot.scala 39:40:@1733.8]
  wire  _T_218; // @[OneHot.scala 39:40:@1734.8]
  wire  _T_219; // @[OneHot.scala 39:40:@1735.8]
  wire [3:0] _T_237; // @[Mux.scala 31:69:@1737.8]
  wire [3:0] _T_238; // @[Mux.scala 31:69:@1738.8]
  wire [3:0] _T_239; // @[Mux.scala 31:69:@1739.8]
  wire [3:0] _T_240; // @[Mux.scala 31:69:@1740.8]
  wire [3:0] _T_241; // @[Mux.scala 31:69:@1741.8]
  wire [3:0] _T_242; // @[Mux.scala 31:69:@1742.8]
  wire [3:0] _T_243; // @[Mux.scala 31:69:@1743.8]
  wire [3:0] _T_244; // @[Mux.scala 31:69:@1744.8]
  wire [3:0] _T_245; // @[Mux.scala 31:69:@1745.8]
  wire [3:0] _T_246; // @[Mux.scala 31:69:@1746.8]
  wire [3:0] _T_247; // @[Mux.scala 31:69:@1747.8]
  wire [3:0] _T_248; // @[Mux.scala 31:69:@1748.8]
  wire [3:0] _T_249; // @[Mux.scala 31:69:@1749.8]
  wire [3:0] _T_250; // @[Mux.scala 31:69:@1750.8]
  wire [3:0] _T_251; // @[Mux.scala 31:69:@1751.8]
  wire [4:0] _GEN_29; // @[Arithmetic_Logic_Unit.scala 130:38:@1678.6]
  wire [65550:0] _GEN_30; // @[Arithmetic_Logic_Unit.scala 129:65:@1676.4]
  wire  _T_253; // @[Arithmetic_Logic_Unit.scala 136:49:@1755.4]
  wire  _T_257; // @[OneHot.scala 39:40:@1762.8]
  wire  _T_258; // @[OneHot.scala 39:40:@1763.8]
  wire  _T_259; // @[OneHot.scala 39:40:@1764.8]
  wire  _T_260; // @[OneHot.scala 39:40:@1765.8]
  wire  _T_261; // @[OneHot.scala 39:40:@1766.8]
  wire  _T_262; // @[OneHot.scala 39:40:@1767.8]
  wire  _T_263; // @[OneHot.scala 39:40:@1768.8]
  wire  _T_264; // @[OneHot.scala 39:40:@1769.8]
  wire  _T_265; // @[OneHot.scala 39:40:@1770.8]
  wire  _T_266; // @[OneHot.scala 39:40:@1771.8]
  wire  _T_267; // @[OneHot.scala 39:40:@1772.8]
  wire  _T_268; // @[OneHot.scala 39:40:@1773.8]
  wire  _T_269; // @[OneHot.scala 39:40:@1774.8]
  wire  _T_270; // @[OneHot.scala 39:40:@1775.8]
  wire  _T_271; // @[OneHot.scala 39:40:@1776.8]
  wire [3:0] _T_289; // @[Mux.scala 31:69:@1778.8]
  wire [3:0] _T_290; // @[Mux.scala 31:69:@1779.8]
  wire [3:0] _T_291; // @[Mux.scala 31:69:@1780.8]
  wire [3:0] _T_292; // @[Mux.scala 31:69:@1781.8]
  wire [3:0] _T_293; // @[Mux.scala 31:69:@1782.8]
  wire [3:0] _T_294; // @[Mux.scala 31:69:@1783.8]
  wire [3:0] _T_295; // @[Mux.scala 31:69:@1784.8]
  wire [3:0] _T_296; // @[Mux.scala 31:69:@1785.8]
  wire [3:0] _T_297; // @[Mux.scala 31:69:@1786.8]
  wire [3:0] _T_298; // @[Mux.scala 31:69:@1787.8]
  wire [3:0] _T_299; // @[Mux.scala 31:69:@1788.8]
  wire [3:0] _T_300; // @[Mux.scala 31:69:@1789.8]
  wire [3:0] _T_301; // @[Mux.scala 31:69:@1790.8]
  wire [3:0] _T_302; // @[Mux.scala 31:69:@1791.8]
  wire [3:0] _T_303; // @[Mux.scala 31:69:@1792.8]
  wire [4:0] _GEN_31; // @[Arithmetic_Logic_Unit.scala 137:39:@1758.6]
  wire [65550:0] _GEN_32; // @[Arithmetic_Logic_Unit.scala 136:65:@1756.4]
  wire  _T_305; // @[Arithmetic_Logic_Unit.scala 143:50:@1796.4]
  wire [65550:0] _GEN_33; // @[Arithmetic_Logic_Unit.scala 143:67:@1797.4]
  wire  _T_377; // @[Arithmetic_Logic_Unit.scala 171:58:@1834.4]
  wire  _T_378; // @[Arithmetic_Logic_Unit.scala 171:58:@1835.4]
  wire  _T_379; // @[Arithmetic_Logic_Unit.scala 171:58:@1836.4]
  wire  _T_380; // @[Arithmetic_Logic_Unit.scala 171:58:@1837.4]
  wire  _T_381; // @[Arithmetic_Logic_Unit.scala 171:58:@1838.4]
  wire  _T_382; // @[Arithmetic_Logic_Unit.scala 171:58:@1839.4]
  wire  _T_383; // @[Arithmetic_Logic_Unit.scala 171:58:@1840.4]
  wire  _T_384; // @[Arithmetic_Logic_Unit.scala 171:58:@1841.4]
  wire  _T_385; // @[Arithmetic_Logic_Unit.scala 171:58:@1842.4]
  wire  _T_386; // @[Arithmetic_Logic_Unit.scala 171:58:@1843.4]
  wire  _T_387; // @[Arithmetic_Logic_Unit.scala 171:58:@1844.4]
  wire  _T_388; // @[Arithmetic_Logic_Unit.scala 171:58:@1845.4]
  wire  _T_389; // @[Arithmetic_Logic_Unit.scala 171:58:@1846.4]
  wire  _T_390; // @[Arithmetic_Logic_Unit.scala 171:58:@1847.4]
  wire  _T_391; // @[Arithmetic_Logic_Unit.scala 171:58:@1848.4]
  wire  _T_392; // @[Arithmetic_Logic_Unit.scala 171:58:@1849.4]
  wire  _T_393; // @[Arithmetic_Logic_Unit.scala 171:58:@1850.4]
  wire  _T_394; // @[Arithmetic_Logic_Unit.scala 171:58:@1851.4]
  wire  _T_395; // @[Arithmetic_Logic_Unit.scala 171:58:@1852.4]
  wire  _T_396; // @[Arithmetic_Logic_Unit.scala 171:58:@1853.4]
  wire  _T_397; // @[Arithmetic_Logic_Unit.scala 171:58:@1854.4]
  wire  _T_398; // @[Arithmetic_Logic_Unit.scala 171:58:@1855.4]
  wire  _T_399; // @[Arithmetic_Logic_Unit.scala 171:58:@1856.4]
  wire  _T_400; // @[Arithmetic_Logic_Unit.scala 171:58:@1857.4]
  wire  _T_401; // @[Arithmetic_Logic_Unit.scala 171:58:@1858.4]
  wire  _T_402; // @[Arithmetic_Logic_Unit.scala 171:58:@1859.4]
  wire  _T_403; // @[Arithmetic_Logic_Unit.scala 171:58:@1860.4]
  wire  _T_404; // @[Arithmetic_Logic_Unit.scala 171:58:@1861.4]
  wire  _T_405; // @[Arithmetic_Logic_Unit.scala 171:58:@1862.4]
  wire  _T_406; // @[Arithmetic_Logic_Unit.scala 171:58:@1863.4]
  wire  _T_407; // @[Arithmetic_Logic_Unit.scala 171:58:@1864.4]
  wire  _T_410; // @[Arithmetic_Logic_Unit.scala 171:55:@1866.4]
  wire  _T_411; // @[Arithmetic_Logic_Unit.scala 171:55:@1867.4]
  wire  _T_412; // @[Arithmetic_Logic_Unit.scala 171:55:@1868.4]
  wire  _T_413; // @[Arithmetic_Logic_Unit.scala 171:55:@1869.4]
  wire  _T_414; // @[Arithmetic_Logic_Unit.scala 171:55:@1870.4]
  wire  _T_415; // @[Arithmetic_Logic_Unit.scala 171:55:@1871.4]
  wire  _T_416; // @[Arithmetic_Logic_Unit.scala 171:55:@1872.4]
  wire  _T_417; // @[Arithmetic_Logic_Unit.scala 171:55:@1873.4]
  wire  _T_418; // @[Arithmetic_Logic_Unit.scala 171:55:@1874.4]
  wire  _T_419; // @[Arithmetic_Logic_Unit.scala 171:55:@1875.4]
  wire  _T_420; // @[Arithmetic_Logic_Unit.scala 171:55:@1876.4]
  wire  _T_421; // @[Arithmetic_Logic_Unit.scala 171:55:@1877.4]
  wire  _T_422; // @[Arithmetic_Logic_Unit.scala 171:55:@1878.4]
  wire  _T_423; // @[Arithmetic_Logic_Unit.scala 171:55:@1879.4]
  wire  _T_424; // @[Arithmetic_Logic_Unit.scala 171:55:@1880.4]
  wire  _T_425; // @[Arithmetic_Logic_Unit.scala 171:55:@1881.4]
  wire  _T_426; // @[Arithmetic_Logic_Unit.scala 171:55:@1882.4]
  wire  _T_427; // @[Arithmetic_Logic_Unit.scala 171:55:@1883.4]
  wire  _T_428; // @[Arithmetic_Logic_Unit.scala 171:55:@1884.4]
  wire  _T_429; // @[Arithmetic_Logic_Unit.scala 171:55:@1885.4]
  wire  _T_430; // @[Arithmetic_Logic_Unit.scala 171:55:@1886.4]
  wire  _T_431; // @[Arithmetic_Logic_Unit.scala 171:55:@1887.4]
  wire  _T_432; // @[Arithmetic_Logic_Unit.scala 171:55:@1888.4]
  wire  _T_433; // @[Arithmetic_Logic_Unit.scala 171:55:@1889.4]
  wire  _T_434; // @[Arithmetic_Logic_Unit.scala 171:55:@1890.4]
  wire  _T_435; // @[Arithmetic_Logic_Unit.scala 171:55:@1891.4]
  wire  _T_436; // @[Arithmetic_Logic_Unit.scala 171:55:@1892.4]
  wire  _T_437; // @[Arithmetic_Logic_Unit.scala 171:55:@1893.4]
  wire  _T_438; // @[Arithmetic_Logic_Unit.scala 171:55:@1894.4]
  wire  _T_439; // @[Arithmetic_Logic_Unit.scala 171:55:@1895.4]
  wire [15:0] result_unsigned; // @[Arithmetic_Logic_Unit.scala 65:29:@1489.4 Arithmetic_Logic_Unit.scala 66:40:@1491.4 Arithmetic_Logic_Unit.scala 78:19:@1502.4 Arithmetic_Logic_Unit.scala 95:82:@1508.6 Arithmetic_Logic_Unit.scala 96:82:@1512.6 Arithmetic_Logic_Unit.scala 97:82:@1518.6 Arithmetic_Logic_Unit.scala 98:82:@1525.6 Arithmetic_Logic_Unit.scala 99:82:@1531.6 Arithmetic_Logic_Unit.scala 100:82:@1536.6 Arithmetic_Logic_Unit.scala 101:80:@1541.6 Arithmetic_Logic_Unit.scala 102:80:@1546.6 Arithmetic_Logic_Unit.scala 103:82:@1551.6 Arithmetic_Logic_Unit.scala 104:83:@1556.6 Arithmetic_Logic_Unit.scala 105:82:@1561.6 Arithmetic_Logic_Unit.scala 106:82:@1566.6 Arithmetic_Logic_Unit.scala 107:84:@1571.6 Arithmetic_Logic_Unit.scala 108:86:@1577.6 Arithmetic_Logic_Unit.scala 109:82:@1582.6 Arithmetic_Logic_Unit.scala 110:84:@1588.6 Arithmetic_Logic_Unit.scala 111:84:@1593.6 Arithmetic_Logic_Unit.scala 112:86:@1599.6 Arithmetic_Logic_Unit.scala 113:84:@1604.6 Arithmetic_Logic_Unit.scala 114:86:@1610.6 Arithmetic_Logic_Unit.scala 115:82:@1615.6 Arithmetic_Logic_Unit.scala 116:84:@1621.6 Arithmetic_Logic_Unit.scala 117:84:@1628.6 Arithmetic_Logic_Unit.scala 118:86:@1636.6 Arithmetic_Logic_Unit.scala 119:80:@1642.6 Arithmetic_Logic_Unit.scala 122:25:@1650.8 Arithmetic_Logic_Unit.scala 124:25:@1657.8 Arithmetic_Logic_Unit.scala 127:80:@1666.6 Arithmetic_Logic_Unit.scala 128:80:@1673.6 Arithmetic_Logic_Unit.scala 131:25:@1679.8 Arithmetic_Logic_Unit.scala 133:25:@1752.8 Arithmetic_Logic_Unit.scala 138:25:@1759.8 Arithmetic_Logic_Unit.scala 140:25:@1793.8 Arithmetic_Logic_Unit.scala 144:23:@1798.6]
  wire  _T_530; // @[Arithmetic_Logic_Unit.scala 181:9:@1968.4]
  assign logical_operand0_unsigned = io_0 != 16'h0; // @[Arithmetic_Logic_Unit.scala 91:58:@1503.4]
  assign logical_operand1_unsigned = io_1 != 16'h0; // @[Arithmetic_Logic_Unit.scala 92:58:@1504.4]
  assign logical_operand2_unsigned = io_3 != 16'h0; // @[Arithmetic_Logic_Unit.scala 93:58:@1505.4]
  assign _T_43 = io_4 == 5'h1; // @[Arithmetic_Logic_Unit.scala 96:49:@1510.4]
  assign _GEN_1 = _T_43 ? io_0 : 16'h0; // @[Arithmetic_Logic_Unit.scala 96:65:@1511.4]
  assign _T_45 = io_4 == 5'h2; // @[Arithmetic_Logic_Unit.scala 97:49:@1514.4]
  assign _T_46 = io_0 + io_1; // @[Arithmetic_Logic_Unit.scala 97:103:@1516.6]
  assign _T_47 = io_0 + io_1; // @[Arithmetic_Logic_Unit.scala 97:103:@1517.6]
  assign _GEN_2 = _T_45 ? _T_47 : _GEN_1; // @[Arithmetic_Logic_Unit.scala 97:65:@1515.4]
  assign _T_49 = io_4 == 5'h3; // @[Arithmetic_Logic_Unit.scala 98:49:@1520.4]
  assign _T_50 = io_0 - io_1; // @[Arithmetic_Logic_Unit.scala 98:103:@1522.6]
  assign _T_51 = $unsigned(_T_50); // @[Arithmetic_Logic_Unit.scala 98:103:@1523.6]
  assign _T_52 = _T_51[15:0]; // @[Arithmetic_Logic_Unit.scala 98:103:@1524.6]
  assign _GEN_3 = _T_49 ? _T_52 : _GEN_2; // @[Arithmetic_Logic_Unit.scala 98:65:@1521.4]
  assign _T_54 = io_4 == 5'h4; // @[Arithmetic_Logic_Unit.scala 99:49:@1527.4]
  assign _GEN_37 = {{65535'd0}, io_0}; // @[Arithmetic_Logic_Unit.scala 99:103:@1530.6]
  assign _T_56 = _GEN_37 << io_1; // @[Arithmetic_Logic_Unit.scala 99:103:@1530.6]
  assign _GEN_4 = _T_54 ? _T_56 : {{65535'd0}, _GEN_3}; // @[Arithmetic_Logic_Unit.scala 99:65:@1528.4]
  assign _T_58 = io_4 == 5'h6; // @[Arithmetic_Logic_Unit.scala 100:49:@1533.4]
  assign _T_59 = io_0 >> io_1; // @[Arithmetic_Logic_Unit.scala 100:103:@1535.6]
  assign _GEN_5 = _T_58 ? {{65535'd0}, _T_59} : _GEN_4; // @[Arithmetic_Logic_Unit.scala 100:65:@1534.4]
  assign _T_61 = io_4 == 5'h7; // @[Arithmetic_Logic_Unit.scala 101:48:@1538.4]
  assign _T_62 = io_0 == io_1; // @[Arithmetic_Logic_Unit.scala 101:101:@1540.6]
  assign _GEN_6 = _T_61 ? {{65550'd0}, _T_62} : _GEN_5; // @[Arithmetic_Logic_Unit.scala 101:63:@1539.4]
  assign _T_64 = io_4 == 5'h8; // @[Arithmetic_Logic_Unit.scala 102:48:@1543.4]
  assign _T_65 = io_0 != io_1; // @[Arithmetic_Logic_Unit.scala 102:101:@1545.6]
  assign _GEN_7 = _T_64 ? {{65550'd0}, _T_65} : _GEN_6; // @[Arithmetic_Logic_Unit.scala 102:63:@1544.4]
  assign _T_67 = io_4 == 5'ha; // @[Arithmetic_Logic_Unit.scala 103:49:@1548.4]
  assign _T_68 = io_0 > io_1; // @[Arithmetic_Logic_Unit.scala 103:103:@1550.6]
  assign _GEN_8 = _T_67 ? {{65550'd0}, _T_68} : _GEN_7; // @[Arithmetic_Logic_Unit.scala 103:65:@1549.4]
  assign _T_70 = io_4 == 5'hc; // @[Arithmetic_Logic_Unit.scala 104:49:@1553.4]
  assign _T_71 = io_0 < io_1; // @[Arithmetic_Logic_Unit.scala 104:104:@1555.6]
  assign _GEN_9 = _T_70 ? {{65550'd0}, _T_71} : _GEN_8; // @[Arithmetic_Logic_Unit.scala 104:66:@1554.4]
  assign _T_73 = io_4 == 5'he; // @[Arithmetic_Logic_Unit.scala 105:49:@1558.4]
  assign _T_74 = io_0 >= io_1; // @[Arithmetic_Logic_Unit.scala 105:103:@1560.6]
  assign _GEN_10 = _T_73 ? {{65550'd0}, _T_74} : _GEN_9; // @[Arithmetic_Logic_Unit.scala 105:65:@1559.4]
  assign _T_76 = io_4 == 5'h10; // @[Arithmetic_Logic_Unit.scala 106:49:@1563.4]
  assign _T_77 = io_0 <= io_1; // @[Arithmetic_Logic_Unit.scala 106:103:@1565.6]
  assign _GEN_11 = _T_76 ? {{65550'd0}, _T_77} : _GEN_10; // @[Arithmetic_Logic_Unit.scala 106:65:@1564.4]
  assign _T_79 = io_4 == 5'h11; // @[Arithmetic_Logic_Unit.scala 107:50:@1568.4]
  assign _T_80 = io_0 & io_1; // @[Arithmetic_Logic_Unit.scala 107:105:@1570.6]
  assign _GEN_12 = _T_79 ? {{65535'd0}, _T_80} : _GEN_11; // @[Arithmetic_Logic_Unit.scala 107:67:@1569.4]
  assign _T_82 = io_4 == 5'h12; // @[Arithmetic_Logic_Unit.scala 108:51:@1573.4]
  assign _T_84 = ~ _T_80; // @[Arithmetic_Logic_Unit.scala 108:89:@1576.6]
  assign _GEN_13 = _T_82 ? {{65535'd0}, _T_84} : _GEN_12; // @[Arithmetic_Logic_Unit.scala 108:69:@1574.4]
  assign _T_86 = io_4 == 5'h13; // @[Arithmetic_Logic_Unit.scala 109:49:@1579.4]
  assign _T_87 = io_0 | io_1; // @[Arithmetic_Logic_Unit.scala 109:103:@1581.6]
  assign _GEN_14 = _T_86 ? {{65535'd0}, _T_87} : _GEN_13; // @[Arithmetic_Logic_Unit.scala 109:65:@1580.4]
  assign _T_89 = io_4 == 5'h14; // @[Arithmetic_Logic_Unit.scala 110:50:@1584.4]
  assign _T_91 = ~ _T_87; // @[Arithmetic_Logic_Unit.scala 110:87:@1587.6]
  assign _GEN_15 = _T_89 ? {{65535'd0}, _T_91} : _GEN_14; // @[Arithmetic_Logic_Unit.scala 110:67:@1585.4]
  assign _T_93 = io_4 == 5'h15; // @[Arithmetic_Logic_Unit.scala 111:50:@1590.4]
  assign _T_94 = io_0 ^ io_1; // @[Arithmetic_Logic_Unit.scala 111:105:@1592.6]
  assign _GEN_16 = _T_93 ? {{65535'd0}, _T_94} : _GEN_15; // @[Arithmetic_Logic_Unit.scala 111:67:@1591.4]
  assign _T_96 = io_4 == 5'h16; // @[Arithmetic_Logic_Unit.scala 112:51:@1595.4]
  assign _T_98 = ~ _T_94; // @[Arithmetic_Logic_Unit.scala 112:89:@1598.6]
  assign _GEN_17 = _T_96 ? {{65535'd0}, _T_98} : _GEN_16; // @[Arithmetic_Logic_Unit.scala 112:69:@1596.4]
  assign _T_100 = io_4 == 5'h17; // @[Arithmetic_Logic_Unit.scala 113:50:@1601.4]
  assign _T_101 = logical_operand0_unsigned & logical_operand1_unsigned; // @[Arithmetic_Logic_Unit.scala 113:113:@1603.6]
  assign _GEN_18 = _T_100 ? {{65550'd0}, _T_101} : _GEN_17; // @[Arithmetic_Logic_Unit.scala 113:67:@1602.4]
  assign _T_103 = io_4 == 5'h18; // @[Arithmetic_Logic_Unit.scala 114:51:@1606.4]
  assign _T_106 = _T_101 == 1'h0; // @[Arithmetic_Logic_Unit.scala 114:89:@1609.6]
  assign _GEN_19 = _T_103 ? {{65550'd0}, _T_106} : _GEN_18; // @[Arithmetic_Logic_Unit.scala 114:69:@1607.4]
  assign _T_108 = io_4 == 5'h19; // @[Arithmetic_Logic_Unit.scala 115:49:@1612.4]
  assign _T_109 = logical_operand0_unsigned | logical_operand1_unsigned; // @[Arithmetic_Logic_Unit.scala 115:111:@1614.6]
  assign _GEN_20 = _T_108 ? {{65550'd0}, _T_109} : _GEN_19; // @[Arithmetic_Logic_Unit.scala 115:65:@1613.4]
  assign _T_111 = io_4 == 5'h1a; // @[Arithmetic_Logic_Unit.scala 116:50:@1617.4]
  assign _T_114 = _T_109 == 1'h0; // @[Arithmetic_Logic_Unit.scala 116:87:@1620.6]
  assign _GEN_21 = _T_111 ? {{65550'd0}, _T_114} : _GEN_20; // @[Arithmetic_Logic_Unit.scala 116:67:@1618.4]
  assign _T_116 = io_4 == 5'h1b; // @[Arithmetic_Logic_Unit.scala 117:50:@1623.4]
  assign _T_118 = logical_operand0_unsigned == 1'h0; // @[Arithmetic_Logic_Unit.scala 117:87:@1625.6]
  assign _T_120 = logical_operand1_unsigned == 1'h0; // @[Arithmetic_Logic_Unit.scala 117:116:@1626.6]
  assign _T_121 = _T_118 ^ _T_120; // @[Arithmetic_Logic_Unit.scala 117:114:@1627.6]
  assign _GEN_22 = _T_116 ? {{65550'd0}, _T_121} : _GEN_21; // @[Arithmetic_Logic_Unit.scala 117:67:@1624.4]
  assign _T_123 = io_4 == 5'h1c; // @[Arithmetic_Logic_Unit.scala 118:51:@1630.4]
  assign _T_130 = _T_121 == 1'h0; // @[Arithmetic_Logic_Unit.scala 118:89:@1635.6]
  assign _GEN_23 = _T_123 ? {{65550'd0}, _T_130} : _GEN_22; // @[Arithmetic_Logic_Unit.scala 118:69:@1631.4]
  assign _GEN_38 = {{1'd0}, io_4}; // @[Arithmetic_Logic_Unit.scala 119:48:@1638.4]
  assign _T_132 = _GEN_38 == 6'h21; // @[Arithmetic_Logic_Unit.scala 119:48:@1638.4]
  assign _T_134 = _T_59[0]; // @[Arithmetic_Logic_Unit.scala 119:100:@1641.6]
  assign _GEN_24 = _T_132 ? {{65550'd0}, _T_134} : _GEN_23; // @[Arithmetic_Logic_Unit.scala 119:63:@1639.4]
  assign _T_136 = _GEN_38 == 6'h22; // @[Arithmetic_Logic_Unit.scala 120:48:@1644.4]
  assign _T_139 = 65536'h1 << io_1; // @[Arithmetic_Logic_Unit.scala 122:53:@1648.8]
  assign _GEN_40 = {{65520'd0}, io_0}; // @[Arithmetic_Logic_Unit.scala 122:46:@1649.8]
  assign _T_140 = _GEN_40 | _T_139; // @[Arithmetic_Logic_Unit.scala 122:46:@1649.8]
  assign _T_144 = ~ _T_139; // @[Arithmetic_Logic_Unit.scala 124:49:@1655.8]
  assign _T_145 = _GEN_40 & _T_144; // @[Arithmetic_Logic_Unit.scala 124:46:@1656.8]
  assign _GEN_25 = logical_operand2_unsigned ? _T_140 : _T_145; // @[Arithmetic_Logic_Unit.scala 121:38:@1646.6]
  assign _GEN_26 = _T_136 ? {{15'd0}, _GEN_25} : _GEN_24; // @[Arithmetic_Logic_Unit.scala 120:63:@1645.4]
  assign _T_147 = _GEN_38 == 6'h23; // @[Arithmetic_Logic_Unit.scala 127:48:@1660.4]
  assign _GEN_27 = _T_147 ? {{15'd0}, _T_145} : _GEN_26; // @[Arithmetic_Logic_Unit.scala 127:63:@1661.4]
  assign _T_154 = _GEN_38 == 6'h24; // @[Arithmetic_Logic_Unit.scala 128:48:@1668.4]
  assign _GEN_28 = _T_154 ? {{15'd0}, _T_140} : _GEN_27; // @[Arithmetic_Logic_Unit.scala 128:63:@1669.4]
  assign _T_160 = _GEN_38 == 6'h25; // @[Arithmetic_Logic_Unit.scala 129:49:@1675.4]
  assign _T_162 = io_0 == 16'h0; // @[Arithmetic_Logic_Unit.scala 130:30:@1677.6]
  assign _T_168 = io_0[15:8]; // @[Bitwise.scala 103:21:@1684.8]
  assign _T_169 = {{8'd0}, _T_168}; // @[Bitwise.scala 103:31:@1685.8]
  assign _T_170 = io_0[7:0]; // @[Bitwise.scala 103:46:@1686.8]
  assign _GEN_47 = {{8'd0}, _T_170}; // @[Bitwise.scala 103:65:@1687.8]
  assign _T_171 = _GEN_47 << 8; // @[Bitwise.scala 103:65:@1687.8]
  assign _T_173 = _T_171 & 16'hff00; // @[Bitwise.scala 103:75:@1689.8]
  assign _T_174 = _T_169 | _T_173; // @[Bitwise.scala 103:39:@1690.8]
  assign _T_178 = _T_174[15:4]; // @[Bitwise.scala 103:21:@1694.8]
  assign _GEN_48 = {{4'd0}, _T_178}; // @[Bitwise.scala 103:31:@1695.8]
  assign _T_179 = _GEN_48 & 16'hf0f; // @[Bitwise.scala 103:31:@1695.8]
  assign _T_180 = _T_174[11:0]; // @[Bitwise.scala 103:46:@1696.8]
  assign _GEN_49 = {{4'd0}, _T_180}; // @[Bitwise.scala 103:65:@1697.8]
  assign _T_181 = _GEN_49 << 4; // @[Bitwise.scala 103:65:@1697.8]
  assign _T_183 = _T_181 & 16'hf0f0; // @[Bitwise.scala 103:75:@1699.8]
  assign _T_184 = _T_179 | _T_183; // @[Bitwise.scala 103:39:@1700.8]
  assign _T_188 = _T_184[15:2]; // @[Bitwise.scala 103:21:@1704.8]
  assign _GEN_50 = {{2'd0}, _T_188}; // @[Bitwise.scala 103:31:@1705.8]
  assign _T_189 = _GEN_50 & 16'h3333; // @[Bitwise.scala 103:31:@1705.8]
  assign _T_190 = _T_184[13:0]; // @[Bitwise.scala 103:46:@1706.8]
  assign _GEN_51 = {{2'd0}, _T_190}; // @[Bitwise.scala 103:65:@1707.8]
  assign _T_191 = _GEN_51 << 2; // @[Bitwise.scala 103:65:@1707.8]
  assign _T_193 = _T_191 & 16'hcccc; // @[Bitwise.scala 103:75:@1709.8]
  assign _T_194 = _T_189 | _T_193; // @[Bitwise.scala 103:39:@1710.8]
  assign _T_198 = _T_194[15:1]; // @[Bitwise.scala 103:21:@1714.8]
  assign _GEN_52 = {{1'd0}, _T_198}; // @[Bitwise.scala 103:31:@1715.8]
  assign _T_199 = _GEN_52 & 16'h5555; // @[Bitwise.scala 103:31:@1715.8]
  assign _T_200 = _T_194[14:0]; // @[Bitwise.scala 103:46:@1716.8]
  assign _GEN_53 = {{1'd0}, _T_200}; // @[Bitwise.scala 103:65:@1717.8]
  assign _T_201 = _GEN_53 << 1; // @[Bitwise.scala 103:65:@1717.8]
  assign _T_203 = _T_201 & 16'haaaa; // @[Bitwise.scala 103:75:@1719.8]
  assign _T_204 = _T_199 | _T_203; // @[Bitwise.scala 103:39:@1720.8]
  assign _T_205 = _T_204[0]; // @[OneHot.scala 39:40:@1721.8]
  assign _T_206 = _T_204[1]; // @[OneHot.scala 39:40:@1722.8]
  assign _T_207 = _T_204[2]; // @[OneHot.scala 39:40:@1723.8]
  assign _T_208 = _T_204[3]; // @[OneHot.scala 39:40:@1724.8]
  assign _T_209 = _T_204[4]; // @[OneHot.scala 39:40:@1725.8]
  assign _T_210 = _T_204[5]; // @[OneHot.scala 39:40:@1726.8]
  assign _T_211 = _T_204[6]; // @[OneHot.scala 39:40:@1727.8]
  assign _T_212 = _T_204[7]; // @[OneHot.scala 39:40:@1728.8]
  assign _T_213 = _T_204[8]; // @[OneHot.scala 39:40:@1729.8]
  assign _T_214 = _T_204[9]; // @[OneHot.scala 39:40:@1730.8]
  assign _T_215 = _T_204[10]; // @[OneHot.scala 39:40:@1731.8]
  assign _T_216 = _T_204[11]; // @[OneHot.scala 39:40:@1732.8]
  assign _T_217 = _T_204[12]; // @[OneHot.scala 39:40:@1733.8]
  assign _T_218 = _T_204[13]; // @[OneHot.scala 39:40:@1734.8]
  assign _T_219 = _T_204[14]; // @[OneHot.scala 39:40:@1735.8]
  assign _T_237 = _T_219 ? 4'he : 4'hf; // @[Mux.scala 31:69:@1737.8]
  assign _T_238 = _T_218 ? 4'hd : _T_237; // @[Mux.scala 31:69:@1738.8]
  assign _T_239 = _T_217 ? 4'hc : _T_238; // @[Mux.scala 31:69:@1739.8]
  assign _T_240 = _T_216 ? 4'hb : _T_239; // @[Mux.scala 31:69:@1740.8]
  assign _T_241 = _T_215 ? 4'ha : _T_240; // @[Mux.scala 31:69:@1741.8]
  assign _T_242 = _T_214 ? 4'h9 : _T_241; // @[Mux.scala 31:69:@1742.8]
  assign _T_243 = _T_213 ? 4'h8 : _T_242; // @[Mux.scala 31:69:@1743.8]
  assign _T_244 = _T_212 ? 4'h7 : _T_243; // @[Mux.scala 31:69:@1744.8]
  assign _T_245 = _T_211 ? 4'h6 : _T_244; // @[Mux.scala 31:69:@1745.8]
  assign _T_246 = _T_210 ? 4'h5 : _T_245; // @[Mux.scala 31:69:@1746.8]
  assign _T_247 = _T_209 ? 4'h4 : _T_246; // @[Mux.scala 31:69:@1747.8]
  assign _T_248 = _T_208 ? 4'h3 : _T_247; // @[Mux.scala 31:69:@1748.8]
  assign _T_249 = _T_207 ? 4'h2 : _T_248; // @[Mux.scala 31:69:@1749.8]
  assign _T_250 = _T_206 ? 4'h1 : _T_249; // @[Mux.scala 31:69:@1750.8]
  assign _T_251 = _T_205 ? 4'h0 : _T_250; // @[Mux.scala 31:69:@1751.8]
  assign _GEN_29 = _T_162 ? 5'h10 : {{1'd0}, _T_251}; // @[Arithmetic_Logic_Unit.scala 130:38:@1678.6]
  assign _GEN_30 = _T_160 ? {{65546'd0}, _GEN_29} : _GEN_28; // @[Arithmetic_Logic_Unit.scala 129:65:@1676.4]
  assign _T_253 = _GEN_38 == 6'h26; // @[Arithmetic_Logic_Unit.scala 136:49:@1755.4]
  assign _T_257 = io_0[0]; // @[OneHot.scala 39:40:@1762.8]
  assign _T_258 = io_0[1]; // @[OneHot.scala 39:40:@1763.8]
  assign _T_259 = io_0[2]; // @[OneHot.scala 39:40:@1764.8]
  assign _T_260 = io_0[3]; // @[OneHot.scala 39:40:@1765.8]
  assign _T_261 = io_0[4]; // @[OneHot.scala 39:40:@1766.8]
  assign _T_262 = io_0[5]; // @[OneHot.scala 39:40:@1767.8]
  assign _T_263 = io_0[6]; // @[OneHot.scala 39:40:@1768.8]
  assign _T_264 = io_0[7]; // @[OneHot.scala 39:40:@1769.8]
  assign _T_265 = io_0[8]; // @[OneHot.scala 39:40:@1770.8]
  assign _T_266 = io_0[9]; // @[OneHot.scala 39:40:@1771.8]
  assign _T_267 = io_0[10]; // @[OneHot.scala 39:40:@1772.8]
  assign _T_268 = io_0[11]; // @[OneHot.scala 39:40:@1773.8]
  assign _T_269 = io_0[12]; // @[OneHot.scala 39:40:@1774.8]
  assign _T_270 = io_0[13]; // @[OneHot.scala 39:40:@1775.8]
  assign _T_271 = io_0[14]; // @[OneHot.scala 39:40:@1776.8]
  assign _T_289 = _T_271 ? 4'he : 4'hf; // @[Mux.scala 31:69:@1778.8]
  assign _T_290 = _T_270 ? 4'hd : _T_289; // @[Mux.scala 31:69:@1779.8]
  assign _T_291 = _T_269 ? 4'hc : _T_290; // @[Mux.scala 31:69:@1780.8]
  assign _T_292 = _T_268 ? 4'hb : _T_291; // @[Mux.scala 31:69:@1781.8]
  assign _T_293 = _T_267 ? 4'ha : _T_292; // @[Mux.scala 31:69:@1782.8]
  assign _T_294 = _T_266 ? 4'h9 : _T_293; // @[Mux.scala 31:69:@1783.8]
  assign _T_295 = _T_265 ? 4'h8 : _T_294; // @[Mux.scala 31:69:@1784.8]
  assign _T_296 = _T_264 ? 4'h7 : _T_295; // @[Mux.scala 31:69:@1785.8]
  assign _T_297 = _T_263 ? 4'h6 : _T_296; // @[Mux.scala 31:69:@1786.8]
  assign _T_298 = _T_262 ? 4'h5 : _T_297; // @[Mux.scala 31:69:@1787.8]
  assign _T_299 = _T_261 ? 4'h4 : _T_298; // @[Mux.scala 31:69:@1788.8]
  assign _T_300 = _T_260 ? 4'h3 : _T_299; // @[Mux.scala 31:69:@1789.8]
  assign _T_301 = _T_259 ? 4'h2 : _T_300; // @[Mux.scala 31:69:@1790.8]
  assign _T_302 = _T_258 ? 4'h1 : _T_301; // @[Mux.scala 31:69:@1791.8]
  assign _T_303 = _T_257 ? 4'h0 : _T_302; // @[Mux.scala 31:69:@1792.8]
  assign _GEN_31 = _T_162 ? 5'h10 : {{1'd0}, _T_303}; // @[Arithmetic_Logic_Unit.scala 137:39:@1758.6]
  assign _GEN_32 = _T_253 ? {{65546'd0}, _GEN_31} : _GEN_30; // @[Arithmetic_Logic_Unit.scala 136:65:@1756.4]
  assign _T_305 = _GEN_38 == 6'h27; // @[Arithmetic_Logic_Unit.scala 143:50:@1796.4]
  assign _GEN_33 = _T_305 ? 65551'h0 : _GEN_32; // @[Arithmetic_Logic_Unit.scala 143:67:@1797.4]
  assign _T_377 = 6'h0 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1834.4]
  assign _T_378 = 6'h1 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1835.4]
  assign _T_379 = 6'h2 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1836.4]
  assign _T_380 = 6'h3 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1837.4]
  assign _T_381 = 6'h4 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1838.4]
  assign _T_382 = 6'h6 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1839.4]
  assign _T_383 = 6'h7 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1840.4]
  assign _T_384 = 6'h8 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1841.4]
  assign _T_385 = 6'ha == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1842.4]
  assign _T_386 = 6'hc == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1843.4]
  assign _T_387 = 6'he == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1844.4]
  assign _T_388 = 6'h10 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1845.4]
  assign _T_389 = 6'h11 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1846.4]
  assign _T_390 = 6'h12 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1847.4]
  assign _T_391 = 6'h13 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1848.4]
  assign _T_392 = 6'h14 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1849.4]
  assign _T_393 = 6'h15 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1850.4]
  assign _T_394 = 6'h16 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1851.4]
  assign _T_395 = 6'h17 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1852.4]
  assign _T_396 = 6'h18 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1853.4]
  assign _T_397 = 6'h19 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1854.4]
  assign _T_398 = 6'h1a == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1855.4]
  assign _T_399 = 6'h1b == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1856.4]
  assign _T_400 = 6'h1c == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1857.4]
  assign _T_401 = 6'h21 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1858.4]
  assign _T_402 = 6'h22 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1859.4]
  assign _T_403 = 6'h23 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1860.4]
  assign _T_404 = 6'h24 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1861.4]
  assign _T_405 = 6'h25 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1862.4]
  assign _T_406 = 6'h26 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1863.4]
  assign _T_407 = 6'h27 == _GEN_38; // @[Arithmetic_Logic_Unit.scala 171:58:@1864.4]
  assign _T_410 = _T_377 | _T_378; // @[Arithmetic_Logic_Unit.scala 171:55:@1866.4]
  assign _T_411 = _T_410 | _T_379; // @[Arithmetic_Logic_Unit.scala 171:55:@1867.4]
  assign _T_412 = _T_411 | _T_380; // @[Arithmetic_Logic_Unit.scala 171:55:@1868.4]
  assign _T_413 = _T_412 | _T_381; // @[Arithmetic_Logic_Unit.scala 171:55:@1869.4]
  assign _T_414 = _T_413 | _T_382; // @[Arithmetic_Logic_Unit.scala 171:55:@1870.4]
  assign _T_415 = _T_414 | _T_383; // @[Arithmetic_Logic_Unit.scala 171:55:@1871.4]
  assign _T_416 = _T_415 | _T_384; // @[Arithmetic_Logic_Unit.scala 171:55:@1872.4]
  assign _T_417 = _T_416 | _T_385; // @[Arithmetic_Logic_Unit.scala 171:55:@1873.4]
  assign _T_418 = _T_417 | _T_386; // @[Arithmetic_Logic_Unit.scala 171:55:@1874.4]
  assign _T_419 = _T_418 | _T_387; // @[Arithmetic_Logic_Unit.scala 171:55:@1875.4]
  assign _T_420 = _T_419 | _T_388; // @[Arithmetic_Logic_Unit.scala 171:55:@1876.4]
  assign _T_421 = _T_420 | _T_389; // @[Arithmetic_Logic_Unit.scala 171:55:@1877.4]
  assign _T_422 = _T_421 | _T_390; // @[Arithmetic_Logic_Unit.scala 171:55:@1878.4]
  assign _T_423 = _T_422 | _T_391; // @[Arithmetic_Logic_Unit.scala 171:55:@1879.4]
  assign _T_424 = _T_423 | _T_392; // @[Arithmetic_Logic_Unit.scala 171:55:@1880.4]
  assign _T_425 = _T_424 | _T_393; // @[Arithmetic_Logic_Unit.scala 171:55:@1881.4]
  assign _T_426 = _T_425 | _T_394; // @[Arithmetic_Logic_Unit.scala 171:55:@1882.4]
  assign _T_427 = _T_426 | _T_395; // @[Arithmetic_Logic_Unit.scala 171:55:@1883.4]
  assign _T_428 = _T_427 | _T_396; // @[Arithmetic_Logic_Unit.scala 171:55:@1884.4]
  assign _T_429 = _T_428 | _T_397; // @[Arithmetic_Logic_Unit.scala 171:55:@1885.4]
  assign _T_430 = _T_429 | _T_398; // @[Arithmetic_Logic_Unit.scala 171:55:@1886.4]
  assign _T_431 = _T_430 | _T_399; // @[Arithmetic_Logic_Unit.scala 171:55:@1887.4]
  assign _T_432 = _T_431 | _T_400; // @[Arithmetic_Logic_Unit.scala 171:55:@1888.4]
  assign _T_433 = _T_432 | _T_401; // @[Arithmetic_Logic_Unit.scala 171:55:@1889.4]
  assign _T_434 = _T_433 | _T_402; // @[Arithmetic_Logic_Unit.scala 171:55:@1890.4]
  assign _T_435 = _T_434 | _T_403; // @[Arithmetic_Logic_Unit.scala 171:55:@1891.4]
  assign _T_436 = _T_435 | _T_404; // @[Arithmetic_Logic_Unit.scala 171:55:@1892.4]
  assign _T_437 = _T_436 | _T_405; // @[Arithmetic_Logic_Unit.scala 171:55:@1893.4]
  assign _T_438 = _T_437 | _T_406; // @[Arithmetic_Logic_Unit.scala 171:55:@1894.4]
  assign _T_439 = _T_438 | _T_407; // @[Arithmetic_Logic_Unit.scala 171:55:@1895.4]
  assign result_unsigned = _GEN_33[15:0]; // @[Arithmetic_Logic_Unit.scala 65:29:@1489.4 Arithmetic_Logic_Unit.scala 66:40:@1491.4 Arithmetic_Logic_Unit.scala 78:19:@1502.4 Arithmetic_Logic_Unit.scala 95:82:@1508.6 Arithmetic_Logic_Unit.scala 96:82:@1512.6 Arithmetic_Logic_Unit.scala 97:82:@1518.6 Arithmetic_Logic_Unit.scala 98:82:@1525.6 Arithmetic_Logic_Unit.scala 99:82:@1531.6 Arithmetic_Logic_Unit.scala 100:82:@1536.6 Arithmetic_Logic_Unit.scala 101:80:@1541.6 Arithmetic_Logic_Unit.scala 102:80:@1546.6 Arithmetic_Logic_Unit.scala 103:82:@1551.6 Arithmetic_Logic_Unit.scala 104:83:@1556.6 Arithmetic_Logic_Unit.scala 105:82:@1561.6 Arithmetic_Logic_Unit.scala 106:82:@1566.6 Arithmetic_Logic_Unit.scala 107:84:@1571.6 Arithmetic_Logic_Unit.scala 108:86:@1577.6 Arithmetic_Logic_Unit.scala 109:82:@1582.6 Arithmetic_Logic_Unit.scala 110:84:@1588.6 Arithmetic_Logic_Unit.scala 111:84:@1593.6 Arithmetic_Logic_Unit.scala 112:86:@1599.6 Arithmetic_Logic_Unit.scala 113:84:@1604.6 Arithmetic_Logic_Unit.scala 114:86:@1610.6 Arithmetic_Logic_Unit.scala 115:82:@1615.6 Arithmetic_Logic_Unit.scala 116:84:@1621.6 Arithmetic_Logic_Unit.scala 117:84:@1628.6 Arithmetic_Logic_Unit.scala 118:86:@1636.6 Arithmetic_Logic_Unit.scala 119:80:@1642.6 Arithmetic_Logic_Unit.scala 122:25:@1650.8 Arithmetic_Logic_Unit.scala 124:25:@1657.8 Arithmetic_Logic_Unit.scala 127:80:@1666.6 Arithmetic_Logic_Unit.scala 128:80:@1673.6 Arithmetic_Logic_Unit.scala 131:25:@1679.8 Arithmetic_Logic_Unit.scala 133:25:@1752.8 Arithmetic_Logic_Unit.scala 138:25:@1759.8 Arithmetic_Logic_Unit.scala 140:25:@1793.8 Arithmetic_Logic_Unit.scala 144:23:@1798.6]
  assign _T_530 = reset == 1'h0; // @[Arithmetic_Logic_Unit.scala 181:9:@1968.4]
  assign io_2 = _T_439 ? result_unsigned : 16'h0; // @[Arithmetic_Logic_Unit.scala 172:22:@1897.6 Arithmetic_Logic_Unit.scala 174:22:@1918.8 Arithmetic_Logic_Unit.scala 176:22:@1962.10 Arithmetic_Logic_Unit.scala 178:22:@1965.10]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_530) begin
          $fwrite(32'h80000002,"opcode = %d\n",io_4); // @[Arithmetic_Logic_Unit.scala 181:9:@1970.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_530) begin
          $fwrite(32'h80000002,"operand 0 = %d\n",io_0); // @[Arithmetic_Logic_Unit.scala 182:9:@1975.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_530) begin
          $fwrite(32'h80000002,"operand 1 = %d\n",io_1); // @[Arithmetic_Logic_Unit.scala 183:9:@1980.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_530) begin
          $fwrite(32'h80000002,"result = %d\n",io_2); // @[Arithmetic_Logic_Unit.scala 184:9:@1985.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_530) begin
          $fwrite(32'h80000002,"-----------------------------------\n"); // @[Arithmetic_Logic_Unit.scala 185:9:@1990.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Multiplexer_Hw( // @[:@3835.2]
  input  [1:0]  io_4, // @[:@3838.4]
  output [31:0] io_3, // @[:@3838.4]
  input  [31:0] io_2, // @[:@3838.4]
  input  [31:0] io_1, // @[:@3838.4]
  input  [31:0] io_0 // @[:@3838.4]
);
  wire  _T_23; // @[Multiplexer.scala 105:17:@3843.4]
  wire [31:0] _GEN_0; // @[Multiplexer.scala 105:30:@3844.4]
  wire  _T_25; // @[Multiplexer.scala 105:17:@3847.4]
  wire [31:0] _GEN_1; // @[Multiplexer.scala 105:30:@3848.4]
  wire  _T_27; // @[Multiplexer.scala 105:17:@3851.4]
  assign _T_23 = io_4 == 2'h2; // @[Multiplexer.scala 105:17:@3843.4]
  assign _GEN_0 = _T_23 ? io_2 : 32'h0; // @[Multiplexer.scala 105:30:@3844.4]
  assign _T_25 = io_4 == 2'h1; // @[Multiplexer.scala 105:17:@3847.4]
  assign _GEN_1 = _T_25 ? io_1 : _GEN_0; // @[Multiplexer.scala 105:30:@3848.4]
  assign _T_27 = io_4 == 2'h0; // @[Multiplexer.scala 105:17:@3851.4]
  assign io_3 = _T_27 ? io_0 : _GEN_1; // @[Multiplexer.scala 97:9:@3842.4 Multiplexer.scala 106:24:@3845.6 Multiplexer.scala 106:24:@3849.6 Multiplexer.scala 106:24:@3853.6]
endmodule
module Multiplexer_Hw_6( // @[:@3961.2]
  input  [1:0]  io_4, // @[:@3964.4]
  output [15:0] io_3, // @[:@3964.4]
  input  [15:0] io_2, // @[:@3964.4]
  input  [15:0] io_1, // @[:@3964.4]
  input  [15:0] io_0 // @[:@3964.4]
);
  wire  _T_23; // @[Multiplexer.scala 105:17:@3969.4]
  wire [15:0] _GEN_0; // @[Multiplexer.scala 105:30:@3970.4]
  wire  _T_25; // @[Multiplexer.scala 105:17:@3973.4]
  wire [15:0] _GEN_1; // @[Multiplexer.scala 105:30:@3974.4]
  wire  _T_27; // @[Multiplexer.scala 105:17:@3977.4]
  assign _T_23 = io_4 == 2'h2; // @[Multiplexer.scala 105:17:@3969.4]
  assign _GEN_0 = _T_23 ? io_2 : 16'h0; // @[Multiplexer.scala 105:30:@3970.4]
  assign _T_25 = io_4 == 2'h1; // @[Multiplexer.scala 105:17:@3973.4]
  assign _GEN_1 = _T_25 ? io_1 : _GEN_0; // @[Multiplexer.scala 105:30:@3974.4]
  assign _T_27 = io_4 == 2'h0; // @[Multiplexer.scala 105:17:@3977.4]
  assign io_3 = _T_27 ? io_0 : _GEN_1; // @[Multiplexer.scala 97:9:@3968.4 Multiplexer.scala 106:24:@3971.6 Multiplexer.scala 106:24:@3975.6 Multiplexer.scala 106:24:@3979.6]
endmodule
module Dedicated_PE_Hw( // @[:@4213.2]
  input         clock, // @[:@4214.4]
  input         reset, // @[:@4215.4]
  input         io_24_read_req, // @[:@4216.4]
  output        io_24_read_ack, // @[:@4216.4]
  input  [3:0]  io_24_read_index, // @[:@4216.4]
  output [15:0] io_24_read_data, // @[:@4216.4]
  input         io_24_write_req, // @[:@4216.4]
  output        io_24_write_ack, // @[:@4216.4]
  input  [3:0]  io_24_write_index, // @[:@4216.4]
  input  [15:0] io_24_write_data, // @[:@4216.4]
  output [15:0] io_23, // @[:@4216.4]
  output [15:0] io_22, // @[:@4216.4]
  output [15:0] io_21, // @[:@4216.4]
  output [15:0] io_20, // @[:@4216.4]
  output [31:0] io_19, // @[:@4216.4]
  output [31:0] io_18, // @[:@4216.4]
  input  [15:0] io_17, // @[:@4216.4]
  input  [15:0] io_16, // @[:@4216.4]
  input  [15:0] io_15, // @[:@4216.4]
  input  [15:0] io_14, // @[:@4216.4]
  input  [15:0] io_13, // @[:@4216.4]
  input  [15:0] io_12, // @[:@4216.4]
  input  [15:0] io_11, // @[:@4216.4]
  input  [15:0] io_10, // @[:@4216.4]
  input  [15:0] io_9, // @[:@4216.4]
  input  [15:0] io_8, // @[:@4216.4]
  input  [15:0] io_7, // @[:@4216.4]
  input  [15:0] io_6, // @[:@4216.4]
  input  [31:0] io_5, // @[:@4216.4]
  input  [31:0] io_4, // @[:@4216.4]
  input  [31:0] io_3, // @[:@4216.4]
  input  [31:0] io_2, // @[:@4216.4]
  input  [31:0] io_1, // @[:@4216.4]
  input  [31:0] io_0 // @[:@4216.4]
);
  wire  Delay_Pipe_Hw_clock; // @[Dedicated_PE.scala 86:39:@4219.4]
  wire  Delay_Pipe_Hw_reset; // @[Dedicated_PE.scala 86:39:@4219.4]
  wire [2:0] Delay_Pipe_Hw_io_2; // @[Dedicated_PE.scala 86:39:@4219.4]
  wire [31:0] Delay_Pipe_Hw_io_1; // @[Dedicated_PE.scala 86:39:@4219.4]
  wire [31:0] Delay_Pipe_Hw_io_0; // @[Dedicated_PE.scala 86:39:@4219.4]
  wire  Delay_Pipe_Hw_1_clock; // @[Dedicated_PE.scala 86:39:@4222.4]
  wire  Delay_Pipe_Hw_1_reset; // @[Dedicated_PE.scala 86:39:@4222.4]
  wire [1:0] Delay_Pipe_Hw_1_io_2; // @[Dedicated_PE.scala 86:39:@4222.4]
  wire [31:0] Delay_Pipe_Hw_1_io_1; // @[Dedicated_PE.scala 86:39:@4222.4]
  wire [31:0] Delay_Pipe_Hw_1_io_0; // @[Dedicated_PE.scala 86:39:@4222.4]
  wire  Delay_Pipe_Hw_2_clock; // @[Dedicated_PE.scala 86:39:@4225.4]
  wire  Delay_Pipe_Hw_2_reset; // @[Dedicated_PE.scala 86:39:@4225.4]
  wire [1:0] Delay_Pipe_Hw_2_io_2; // @[Dedicated_PE.scala 86:39:@4225.4]
  wire [31:0] Delay_Pipe_Hw_2_io_1; // @[Dedicated_PE.scala 86:39:@4225.4]
  wire [31:0] Delay_Pipe_Hw_2_io_0; // @[Dedicated_PE.scala 86:39:@4225.4]
  wire  Arithmetic_Logic_Unit_Hw_clock; // @[Dedicated_PE.scala 85:32:@4228.4]
  wire  Arithmetic_Logic_Unit_Hw_reset; // @[Dedicated_PE.scala 85:32:@4228.4]
  wire [4:0] Arithmetic_Logic_Unit_Hw_io_4; // @[Dedicated_PE.scala 85:32:@4228.4]
  wire [31:0] Arithmetic_Logic_Unit_Hw_io_3; // @[Dedicated_PE.scala 85:32:@4228.4]
  wire [31:0] Arithmetic_Logic_Unit_Hw_io_2; // @[Dedicated_PE.scala 85:32:@4228.4]
  wire [31:0] Arithmetic_Logic_Unit_Hw_io_1; // @[Dedicated_PE.scala 85:32:@4228.4]
  wire [31:0] Arithmetic_Logic_Unit_Hw_io_0; // @[Dedicated_PE.scala 85:32:@4228.4]
  wire  Delay_Pipe_Hw_3_clock; // @[Dedicated_PE.scala 86:39:@4231.4]
  wire  Delay_Pipe_Hw_3_reset; // @[Dedicated_PE.scala 86:39:@4231.4]
  wire [2:0] Delay_Pipe_Hw_3_io_2; // @[Dedicated_PE.scala 86:39:@4231.4]
  wire [31:0] Delay_Pipe_Hw_3_io_1; // @[Dedicated_PE.scala 86:39:@4231.4]
  wire [31:0] Delay_Pipe_Hw_3_io_0; // @[Dedicated_PE.scala 86:39:@4231.4]
  wire  Delay_Pipe_Hw_4_clock; // @[Dedicated_PE.scala 86:39:@4234.4]
  wire  Delay_Pipe_Hw_4_reset; // @[Dedicated_PE.scala 86:39:@4234.4]
  wire [1:0] Delay_Pipe_Hw_4_io_2; // @[Dedicated_PE.scala 86:39:@4234.4]
  wire [31:0] Delay_Pipe_Hw_4_io_1; // @[Dedicated_PE.scala 86:39:@4234.4]
  wire [31:0] Delay_Pipe_Hw_4_io_0; // @[Dedicated_PE.scala 86:39:@4234.4]
  wire  Delay_Pipe_Hw_5_clock; // @[Dedicated_PE.scala 86:39:@4237.4]
  wire  Delay_Pipe_Hw_5_reset; // @[Dedicated_PE.scala 86:39:@4237.4]
  wire [1:0] Delay_Pipe_Hw_5_io_2; // @[Dedicated_PE.scala 86:39:@4237.4]
  wire [31:0] Delay_Pipe_Hw_5_io_1; // @[Dedicated_PE.scala 86:39:@4237.4]
  wire [31:0] Delay_Pipe_Hw_5_io_0; // @[Dedicated_PE.scala 86:39:@4237.4]
  wire  Arithmetic_Logic_Unit_Hw_1_clock; // @[Dedicated_PE.scala 85:32:@4240.4]
  wire  Arithmetic_Logic_Unit_Hw_1_reset; // @[Dedicated_PE.scala 85:32:@4240.4]
  wire [4:0] Arithmetic_Logic_Unit_Hw_1_io_4; // @[Dedicated_PE.scala 85:32:@4240.4]
  wire [31:0] Arithmetic_Logic_Unit_Hw_1_io_3; // @[Dedicated_PE.scala 85:32:@4240.4]
  wire [31:0] Arithmetic_Logic_Unit_Hw_1_io_2; // @[Dedicated_PE.scala 85:32:@4240.4]
  wire [31:0] Arithmetic_Logic_Unit_Hw_1_io_1; // @[Dedicated_PE.scala 85:32:@4240.4]
  wire [31:0] Arithmetic_Logic_Unit_Hw_1_io_0; // @[Dedicated_PE.scala 85:32:@4240.4]
  wire  Delay_Pipe_Hw_6_clock; // @[Dedicated_PE.scala 86:39:@4243.4]
  wire  Delay_Pipe_Hw_6_reset; // @[Dedicated_PE.scala 86:39:@4243.4]
  wire [2:0] Delay_Pipe_Hw_6_io_2; // @[Dedicated_PE.scala 86:39:@4243.4]
  wire [15:0] Delay_Pipe_Hw_6_io_1; // @[Dedicated_PE.scala 86:39:@4243.4]
  wire [15:0] Delay_Pipe_Hw_6_io_0; // @[Dedicated_PE.scala 86:39:@4243.4]
  wire  Delay_Pipe_Hw_7_clock; // @[Dedicated_PE.scala 86:39:@4246.4]
  wire  Delay_Pipe_Hw_7_reset; // @[Dedicated_PE.scala 86:39:@4246.4]
  wire [1:0] Delay_Pipe_Hw_7_io_2; // @[Dedicated_PE.scala 86:39:@4246.4]
  wire [15:0] Delay_Pipe_Hw_7_io_1; // @[Dedicated_PE.scala 86:39:@4246.4]
  wire [15:0] Delay_Pipe_Hw_7_io_0; // @[Dedicated_PE.scala 86:39:@4246.4]
  wire  Delay_Pipe_Hw_8_clock; // @[Dedicated_PE.scala 86:39:@4249.4]
  wire  Delay_Pipe_Hw_8_reset; // @[Dedicated_PE.scala 86:39:@4249.4]
  wire [1:0] Delay_Pipe_Hw_8_io_2; // @[Dedicated_PE.scala 86:39:@4249.4]
  wire [15:0] Delay_Pipe_Hw_8_io_1; // @[Dedicated_PE.scala 86:39:@4249.4]
  wire [15:0] Delay_Pipe_Hw_8_io_0; // @[Dedicated_PE.scala 86:39:@4249.4]
  wire  Arithmetic_Logic_Unit_Hw_2_clock; // @[Dedicated_PE.scala 85:32:@4252.4]
  wire  Arithmetic_Logic_Unit_Hw_2_reset; // @[Dedicated_PE.scala 85:32:@4252.4]
  wire [4:0] Arithmetic_Logic_Unit_Hw_2_io_4; // @[Dedicated_PE.scala 85:32:@4252.4]
  wire [15:0] Arithmetic_Logic_Unit_Hw_2_io_3; // @[Dedicated_PE.scala 85:32:@4252.4]
  wire [15:0] Arithmetic_Logic_Unit_Hw_2_io_2; // @[Dedicated_PE.scala 85:32:@4252.4]
  wire [15:0] Arithmetic_Logic_Unit_Hw_2_io_1; // @[Dedicated_PE.scala 85:32:@4252.4]
  wire [15:0] Arithmetic_Logic_Unit_Hw_2_io_0; // @[Dedicated_PE.scala 85:32:@4252.4]
  wire  Delay_Pipe_Hw_9_clock; // @[Dedicated_PE.scala 86:39:@4255.4]
  wire  Delay_Pipe_Hw_9_reset; // @[Dedicated_PE.scala 86:39:@4255.4]
  wire [2:0] Delay_Pipe_Hw_9_io_2; // @[Dedicated_PE.scala 86:39:@4255.4]
  wire [15:0] Delay_Pipe_Hw_9_io_1; // @[Dedicated_PE.scala 86:39:@4255.4]
  wire [15:0] Delay_Pipe_Hw_9_io_0; // @[Dedicated_PE.scala 86:39:@4255.4]
  wire  Delay_Pipe_Hw_10_clock; // @[Dedicated_PE.scala 86:39:@4258.4]
  wire  Delay_Pipe_Hw_10_reset; // @[Dedicated_PE.scala 86:39:@4258.4]
  wire [1:0] Delay_Pipe_Hw_10_io_2; // @[Dedicated_PE.scala 86:39:@4258.4]
  wire [15:0] Delay_Pipe_Hw_10_io_1; // @[Dedicated_PE.scala 86:39:@4258.4]
  wire [15:0] Delay_Pipe_Hw_10_io_0; // @[Dedicated_PE.scala 86:39:@4258.4]
  wire  Delay_Pipe_Hw_11_clock; // @[Dedicated_PE.scala 86:39:@4261.4]
  wire  Delay_Pipe_Hw_11_reset; // @[Dedicated_PE.scala 86:39:@4261.4]
  wire [1:0] Delay_Pipe_Hw_11_io_2; // @[Dedicated_PE.scala 86:39:@4261.4]
  wire [15:0] Delay_Pipe_Hw_11_io_1; // @[Dedicated_PE.scala 86:39:@4261.4]
  wire [15:0] Delay_Pipe_Hw_11_io_0; // @[Dedicated_PE.scala 86:39:@4261.4]
  wire  Arithmetic_Logic_Unit_Hw_3_clock; // @[Dedicated_PE.scala 85:32:@4264.4]
  wire  Arithmetic_Logic_Unit_Hw_3_reset; // @[Dedicated_PE.scala 85:32:@4264.4]
  wire [4:0] Arithmetic_Logic_Unit_Hw_3_io_4; // @[Dedicated_PE.scala 85:32:@4264.4]
  wire [15:0] Arithmetic_Logic_Unit_Hw_3_io_3; // @[Dedicated_PE.scala 85:32:@4264.4]
  wire [15:0] Arithmetic_Logic_Unit_Hw_3_io_2; // @[Dedicated_PE.scala 85:32:@4264.4]
  wire [15:0] Arithmetic_Logic_Unit_Hw_3_io_1; // @[Dedicated_PE.scala 85:32:@4264.4]
  wire [15:0] Arithmetic_Logic_Unit_Hw_3_io_0; // @[Dedicated_PE.scala 85:32:@4264.4]
  wire  Delay_Pipe_Hw_12_clock; // @[Dedicated_PE.scala 86:39:@4267.4]
  wire  Delay_Pipe_Hw_12_reset; // @[Dedicated_PE.scala 86:39:@4267.4]
  wire [2:0] Delay_Pipe_Hw_12_io_2; // @[Dedicated_PE.scala 86:39:@4267.4]
  wire [15:0] Delay_Pipe_Hw_12_io_1; // @[Dedicated_PE.scala 86:39:@4267.4]
  wire [15:0] Delay_Pipe_Hw_12_io_0; // @[Dedicated_PE.scala 86:39:@4267.4]
  wire  Delay_Pipe_Hw_13_clock; // @[Dedicated_PE.scala 86:39:@4270.4]
  wire  Delay_Pipe_Hw_13_reset; // @[Dedicated_PE.scala 86:39:@4270.4]
  wire [1:0] Delay_Pipe_Hw_13_io_2; // @[Dedicated_PE.scala 86:39:@4270.4]
  wire [15:0] Delay_Pipe_Hw_13_io_1; // @[Dedicated_PE.scala 86:39:@4270.4]
  wire [15:0] Delay_Pipe_Hw_13_io_0; // @[Dedicated_PE.scala 86:39:@4270.4]
  wire  Delay_Pipe_Hw_14_clock; // @[Dedicated_PE.scala 86:39:@4273.4]
  wire  Delay_Pipe_Hw_14_reset; // @[Dedicated_PE.scala 86:39:@4273.4]
  wire [1:0] Delay_Pipe_Hw_14_io_2; // @[Dedicated_PE.scala 86:39:@4273.4]
  wire [15:0] Delay_Pipe_Hw_14_io_1; // @[Dedicated_PE.scala 86:39:@4273.4]
  wire [15:0] Delay_Pipe_Hw_14_io_0; // @[Dedicated_PE.scala 86:39:@4273.4]
  wire  Arithmetic_Logic_Unit_Hw_4_clock; // @[Dedicated_PE.scala 85:32:@4276.4]
  wire  Arithmetic_Logic_Unit_Hw_4_reset; // @[Dedicated_PE.scala 85:32:@4276.4]
  wire [4:0] Arithmetic_Logic_Unit_Hw_4_io_4; // @[Dedicated_PE.scala 85:32:@4276.4]
  wire [15:0] Arithmetic_Logic_Unit_Hw_4_io_3; // @[Dedicated_PE.scala 85:32:@4276.4]
  wire [15:0] Arithmetic_Logic_Unit_Hw_4_io_2; // @[Dedicated_PE.scala 85:32:@4276.4]
  wire [15:0] Arithmetic_Logic_Unit_Hw_4_io_1; // @[Dedicated_PE.scala 85:32:@4276.4]
  wire [15:0] Arithmetic_Logic_Unit_Hw_4_io_0; // @[Dedicated_PE.scala 85:32:@4276.4]
  wire  Delay_Pipe_Hw_15_clock; // @[Dedicated_PE.scala 86:39:@4279.4]
  wire  Delay_Pipe_Hw_15_reset; // @[Dedicated_PE.scala 86:39:@4279.4]
  wire [2:0] Delay_Pipe_Hw_15_io_2; // @[Dedicated_PE.scala 86:39:@4279.4]
  wire [15:0] Delay_Pipe_Hw_15_io_1; // @[Dedicated_PE.scala 86:39:@4279.4]
  wire [15:0] Delay_Pipe_Hw_15_io_0; // @[Dedicated_PE.scala 86:39:@4279.4]
  wire  Delay_Pipe_Hw_16_clock; // @[Dedicated_PE.scala 86:39:@4282.4]
  wire  Delay_Pipe_Hw_16_reset; // @[Dedicated_PE.scala 86:39:@4282.4]
  wire [1:0] Delay_Pipe_Hw_16_io_2; // @[Dedicated_PE.scala 86:39:@4282.4]
  wire [15:0] Delay_Pipe_Hw_16_io_1; // @[Dedicated_PE.scala 86:39:@4282.4]
  wire [15:0] Delay_Pipe_Hw_16_io_0; // @[Dedicated_PE.scala 86:39:@4282.4]
  wire  Delay_Pipe_Hw_17_clock; // @[Dedicated_PE.scala 86:39:@4285.4]
  wire  Delay_Pipe_Hw_17_reset; // @[Dedicated_PE.scala 86:39:@4285.4]
  wire [1:0] Delay_Pipe_Hw_17_io_2; // @[Dedicated_PE.scala 86:39:@4285.4]
  wire [15:0] Delay_Pipe_Hw_17_io_1; // @[Dedicated_PE.scala 86:39:@4285.4]
  wire [15:0] Delay_Pipe_Hw_17_io_0; // @[Dedicated_PE.scala 86:39:@4285.4]
  wire  Arithmetic_Logic_Unit_Hw_5_clock; // @[Dedicated_PE.scala 85:32:@4288.4]
  wire  Arithmetic_Logic_Unit_Hw_5_reset; // @[Dedicated_PE.scala 85:32:@4288.4]
  wire [4:0] Arithmetic_Logic_Unit_Hw_5_io_4; // @[Dedicated_PE.scala 85:32:@4288.4]
  wire [15:0] Arithmetic_Logic_Unit_Hw_5_io_3; // @[Dedicated_PE.scala 85:32:@4288.4]
  wire [15:0] Arithmetic_Logic_Unit_Hw_5_io_2; // @[Dedicated_PE.scala 85:32:@4288.4]
  wire [15:0] Arithmetic_Logic_Unit_Hw_5_io_1; // @[Dedicated_PE.scala 85:32:@4288.4]
  wire [15:0] Arithmetic_Logic_Unit_Hw_5_io_0; // @[Dedicated_PE.scala 85:32:@4288.4]
  wire [1:0] Multiplexer_Hw_io_4; // @[Dedicated_PE.scala 84:32:@4291.4]
  wire [31:0] Multiplexer_Hw_io_3; // @[Dedicated_PE.scala 84:32:@4291.4]
  wire [31:0] Multiplexer_Hw_io_2; // @[Dedicated_PE.scala 84:32:@4291.4]
  wire [31:0] Multiplexer_Hw_io_1; // @[Dedicated_PE.scala 84:32:@4291.4]
  wire [31:0] Multiplexer_Hw_io_0; // @[Dedicated_PE.scala 84:32:@4291.4]
  wire [1:0] Multiplexer_Hw_1_io_4; // @[Dedicated_PE.scala 84:32:@4294.4]
  wire [31:0] Multiplexer_Hw_1_io_3; // @[Dedicated_PE.scala 84:32:@4294.4]
  wire [31:0] Multiplexer_Hw_1_io_2; // @[Dedicated_PE.scala 84:32:@4294.4]
  wire [31:0] Multiplexer_Hw_1_io_1; // @[Dedicated_PE.scala 84:32:@4294.4]
  wire [31:0] Multiplexer_Hw_1_io_0; // @[Dedicated_PE.scala 84:32:@4294.4]
  wire [1:0] Multiplexer_Hw_2_io_4; // @[Dedicated_PE.scala 84:32:@4297.4]
  wire [31:0] Multiplexer_Hw_2_io_3; // @[Dedicated_PE.scala 84:32:@4297.4]
  wire [31:0] Multiplexer_Hw_2_io_2; // @[Dedicated_PE.scala 84:32:@4297.4]
  wire [31:0] Multiplexer_Hw_2_io_1; // @[Dedicated_PE.scala 84:32:@4297.4]
  wire [31:0] Multiplexer_Hw_2_io_0; // @[Dedicated_PE.scala 84:32:@4297.4]
  wire [1:0] Multiplexer_Hw_3_io_4; // @[Dedicated_PE.scala 84:32:@4300.4]
  wire [31:0] Multiplexer_Hw_3_io_3; // @[Dedicated_PE.scala 84:32:@4300.4]
  wire [31:0] Multiplexer_Hw_3_io_2; // @[Dedicated_PE.scala 84:32:@4300.4]
  wire [31:0] Multiplexer_Hw_3_io_1; // @[Dedicated_PE.scala 84:32:@4300.4]
  wire [31:0] Multiplexer_Hw_3_io_0; // @[Dedicated_PE.scala 84:32:@4300.4]
  wire [1:0] Multiplexer_Hw_4_io_4; // @[Dedicated_PE.scala 84:32:@4303.4]
  wire [31:0] Multiplexer_Hw_4_io_3; // @[Dedicated_PE.scala 84:32:@4303.4]
  wire [31:0] Multiplexer_Hw_4_io_2; // @[Dedicated_PE.scala 84:32:@4303.4]
  wire [31:0] Multiplexer_Hw_4_io_1; // @[Dedicated_PE.scala 84:32:@4303.4]
  wire [31:0] Multiplexer_Hw_4_io_0; // @[Dedicated_PE.scala 84:32:@4303.4]
  wire [1:0] Multiplexer_Hw_5_io_4; // @[Dedicated_PE.scala 84:32:@4306.4]
  wire [31:0] Multiplexer_Hw_5_io_3; // @[Dedicated_PE.scala 84:32:@4306.4]
  wire [31:0] Multiplexer_Hw_5_io_2; // @[Dedicated_PE.scala 84:32:@4306.4]
  wire [31:0] Multiplexer_Hw_5_io_1; // @[Dedicated_PE.scala 84:32:@4306.4]
  wire [31:0] Multiplexer_Hw_5_io_0; // @[Dedicated_PE.scala 84:32:@4306.4]
  wire [1:0] Multiplexer_Hw_6_io_4; // @[Dedicated_PE.scala 84:32:@4309.4]
  wire [15:0] Multiplexer_Hw_6_io_3; // @[Dedicated_PE.scala 84:32:@4309.4]
  wire [15:0] Multiplexer_Hw_6_io_2; // @[Dedicated_PE.scala 84:32:@4309.4]
  wire [15:0] Multiplexer_Hw_6_io_1; // @[Dedicated_PE.scala 84:32:@4309.4]
  wire [15:0] Multiplexer_Hw_6_io_0; // @[Dedicated_PE.scala 84:32:@4309.4]
  wire [1:0] Multiplexer_Hw_7_io_4; // @[Dedicated_PE.scala 84:32:@4312.4]
  wire [15:0] Multiplexer_Hw_7_io_3; // @[Dedicated_PE.scala 84:32:@4312.4]
  wire [15:0] Multiplexer_Hw_7_io_2; // @[Dedicated_PE.scala 84:32:@4312.4]
  wire [15:0] Multiplexer_Hw_7_io_1; // @[Dedicated_PE.scala 84:32:@4312.4]
  wire [15:0] Multiplexer_Hw_7_io_0; // @[Dedicated_PE.scala 84:32:@4312.4]
  wire [1:0] Multiplexer_Hw_8_io_4; // @[Dedicated_PE.scala 84:32:@4315.4]
  wire [15:0] Multiplexer_Hw_8_io_3; // @[Dedicated_PE.scala 84:32:@4315.4]
  wire [15:0] Multiplexer_Hw_8_io_2; // @[Dedicated_PE.scala 84:32:@4315.4]
  wire [15:0] Multiplexer_Hw_8_io_1; // @[Dedicated_PE.scala 84:32:@4315.4]
  wire [15:0] Multiplexer_Hw_8_io_0; // @[Dedicated_PE.scala 84:32:@4315.4]
  wire [1:0] Multiplexer_Hw_9_io_4; // @[Dedicated_PE.scala 84:32:@4318.4]
  wire [15:0] Multiplexer_Hw_9_io_3; // @[Dedicated_PE.scala 84:32:@4318.4]
  wire [15:0] Multiplexer_Hw_9_io_2; // @[Dedicated_PE.scala 84:32:@4318.4]
  wire [15:0] Multiplexer_Hw_9_io_1; // @[Dedicated_PE.scala 84:32:@4318.4]
  wire [15:0] Multiplexer_Hw_9_io_0; // @[Dedicated_PE.scala 84:32:@4318.4]
  wire [1:0] Multiplexer_Hw_10_io_4; // @[Dedicated_PE.scala 84:32:@4321.4]
  wire [15:0] Multiplexer_Hw_10_io_3; // @[Dedicated_PE.scala 84:32:@4321.4]
  wire [15:0] Multiplexer_Hw_10_io_2; // @[Dedicated_PE.scala 84:32:@4321.4]
  wire [15:0] Multiplexer_Hw_10_io_1; // @[Dedicated_PE.scala 84:32:@4321.4]
  wire [15:0] Multiplexer_Hw_10_io_0; // @[Dedicated_PE.scala 84:32:@4321.4]
  wire [1:0] Multiplexer_Hw_11_io_4; // @[Dedicated_PE.scala 84:32:@4324.4]
  wire [15:0] Multiplexer_Hw_11_io_3; // @[Dedicated_PE.scala 84:32:@4324.4]
  wire [15:0] Multiplexer_Hw_11_io_2; // @[Dedicated_PE.scala 84:32:@4324.4]
  wire [15:0] Multiplexer_Hw_11_io_1; // @[Dedicated_PE.scala 84:32:@4324.4]
  wire [15:0] Multiplexer_Hw_11_io_0; // @[Dedicated_PE.scala 84:32:@4324.4]
  wire [1:0] Multiplexer_Hw_12_io_4; // @[Dedicated_PE.scala 84:32:@4327.4]
  wire [15:0] Multiplexer_Hw_12_io_3; // @[Dedicated_PE.scala 84:32:@4327.4]
  wire [15:0] Multiplexer_Hw_12_io_2; // @[Dedicated_PE.scala 84:32:@4327.4]
  wire [15:0] Multiplexer_Hw_12_io_1; // @[Dedicated_PE.scala 84:32:@4327.4]
  wire [15:0] Multiplexer_Hw_12_io_0; // @[Dedicated_PE.scala 84:32:@4327.4]
  wire [1:0] Multiplexer_Hw_13_io_4; // @[Dedicated_PE.scala 84:32:@4330.4]
  wire [15:0] Multiplexer_Hw_13_io_3; // @[Dedicated_PE.scala 84:32:@4330.4]
  wire [15:0] Multiplexer_Hw_13_io_2; // @[Dedicated_PE.scala 84:32:@4330.4]
  wire [15:0] Multiplexer_Hw_13_io_1; // @[Dedicated_PE.scala 84:32:@4330.4]
  wire [15:0] Multiplexer_Hw_13_io_0; // @[Dedicated_PE.scala 84:32:@4330.4]
  wire [1:0] Multiplexer_Hw_14_io_4; // @[Dedicated_PE.scala 84:32:@4333.4]
  wire [15:0] Multiplexer_Hw_14_io_3; // @[Dedicated_PE.scala 84:32:@4333.4]
  wire [15:0] Multiplexer_Hw_14_io_2; // @[Dedicated_PE.scala 84:32:@4333.4]
  wire [15:0] Multiplexer_Hw_14_io_1; // @[Dedicated_PE.scala 84:32:@4333.4]
  wire [15:0] Multiplexer_Hw_14_io_0; // @[Dedicated_PE.scala 84:32:@4333.4]
  wire [1:0] Multiplexer_Hw_15_io_4; // @[Dedicated_PE.scala 84:32:@4336.4]
  wire [15:0] Multiplexer_Hw_15_io_3; // @[Dedicated_PE.scala 84:32:@4336.4]
  wire [15:0] Multiplexer_Hw_15_io_2; // @[Dedicated_PE.scala 84:32:@4336.4]
  wire [15:0] Multiplexer_Hw_15_io_1; // @[Dedicated_PE.scala 84:32:@4336.4]
  wire [15:0] Multiplexer_Hw_15_io_0; // @[Dedicated_PE.scala 84:32:@4336.4]
  wire [1:0] Multiplexer_Hw_16_io_4; // @[Dedicated_PE.scala 84:32:@4339.4]
  wire [15:0] Multiplexer_Hw_16_io_3; // @[Dedicated_PE.scala 84:32:@4339.4]
  wire [15:0] Multiplexer_Hw_16_io_2; // @[Dedicated_PE.scala 84:32:@4339.4]
  wire [15:0] Multiplexer_Hw_16_io_1; // @[Dedicated_PE.scala 84:32:@4339.4]
  wire [15:0] Multiplexer_Hw_16_io_0; // @[Dedicated_PE.scala 84:32:@4339.4]
  wire [1:0] Multiplexer_Hw_17_io_4; // @[Dedicated_PE.scala 84:32:@4342.4]
  wire [15:0] Multiplexer_Hw_17_io_3; // @[Dedicated_PE.scala 84:32:@4342.4]
  wire [15:0] Multiplexer_Hw_17_io_2; // @[Dedicated_PE.scala 84:32:@4342.4]
  wire [15:0] Multiplexer_Hw_17_io_1; // @[Dedicated_PE.scala 84:32:@4342.4]
  wire [15:0] Multiplexer_Hw_17_io_0; // @[Dedicated_PE.scala 84:32:@4342.4]
  reg [15:0] config_registers_0; // @[Dedicated_PE.scala 76:29:@4218.4]
  reg [31:0] _RAND_0;
  reg [15:0] config_registers_1; // @[Dedicated_PE.scala 76:29:@4218.4]
  reg [31:0] _RAND_1;
  reg [15:0] config_registers_2; // @[Dedicated_PE.scala 76:29:@4218.4]
  reg [31:0] _RAND_2;
  reg [15:0] config_registers_3; // @[Dedicated_PE.scala 76:29:@4218.4]
  reg [31:0] _RAND_3;
  reg [15:0] config_registers_4; // @[Dedicated_PE.scala 76:29:@4218.4]
  reg [31:0] _RAND_4;
  reg [15:0] config_registers_5; // @[Dedicated_PE.scala 76:29:@4218.4]
  reg [31:0] _RAND_5;
  reg [15:0] config_registers_6; // @[Dedicated_PE.scala 76:29:@4218.4]
  reg [31:0] _RAND_6;
  reg [15:0] config_registers_7; // @[Dedicated_PE.scala 76:29:@4218.4]
  reg [31:0] _RAND_7;
  wire [2:0] _T_167; // @[:@4526.6]
  wire [15:0] _GEN_0; // @[Dedicated_PE.scala 137:47:@4527.6]
  wire [15:0] _GEN_1; // @[Dedicated_PE.scala 137:47:@4527.6]
  wire [15:0] _GEN_2; // @[Dedicated_PE.scala 137:47:@4527.6]
  wire [15:0] _GEN_3; // @[Dedicated_PE.scala 137:47:@4527.6]
  wire [15:0] _GEN_4; // @[Dedicated_PE.scala 137:47:@4527.6]
  wire [15:0] _GEN_5; // @[Dedicated_PE.scala 137:47:@4527.6]
  wire [15:0] _GEN_6; // @[Dedicated_PE.scala 137:47:@4527.6]
  wire [15:0] _GEN_7; // @[Dedicated_PE.scala 137:47:@4527.6]
  Delay_Pipe_Hw Delay_Pipe_Hw ( // @[Dedicated_PE.scala 86:39:@4219.4]
    .clock(Delay_Pipe_Hw_clock),
    .reset(Delay_Pipe_Hw_reset),
    .io_2(Delay_Pipe_Hw_io_2),
    .io_1(Delay_Pipe_Hw_io_1),
    .io_0(Delay_Pipe_Hw_io_0)
  );
  Delay_Pipe_Hw_1 Delay_Pipe_Hw_1 ( // @[Dedicated_PE.scala 86:39:@4222.4]
    .clock(Delay_Pipe_Hw_1_clock),
    .reset(Delay_Pipe_Hw_1_reset),
    .io_2(Delay_Pipe_Hw_1_io_2),
    .io_1(Delay_Pipe_Hw_1_io_1),
    .io_0(Delay_Pipe_Hw_1_io_0)
  );
  Delay_Pipe_Hw_1 Delay_Pipe_Hw_2 ( // @[Dedicated_PE.scala 86:39:@4225.4]
    .clock(Delay_Pipe_Hw_2_clock),
    .reset(Delay_Pipe_Hw_2_reset),
    .io_2(Delay_Pipe_Hw_2_io_2),
    .io_1(Delay_Pipe_Hw_2_io_1),
    .io_0(Delay_Pipe_Hw_2_io_0)
  );
  Arithmetic_Logic_Unit_Hw Arithmetic_Logic_Unit_Hw ( // @[Dedicated_PE.scala 85:32:@4228.4]
    .clock(Arithmetic_Logic_Unit_Hw_clock),
    .reset(Arithmetic_Logic_Unit_Hw_reset),
    .io_4(Arithmetic_Logic_Unit_Hw_io_4),
    .io_3(Arithmetic_Logic_Unit_Hw_io_3),
    .io_2(Arithmetic_Logic_Unit_Hw_io_2),
    .io_1(Arithmetic_Logic_Unit_Hw_io_1),
    .io_0(Arithmetic_Logic_Unit_Hw_io_0)
  );
  Delay_Pipe_Hw Delay_Pipe_Hw_3 ( // @[Dedicated_PE.scala 86:39:@4231.4]
    .clock(Delay_Pipe_Hw_3_clock),
    .reset(Delay_Pipe_Hw_3_reset),
    .io_2(Delay_Pipe_Hw_3_io_2),
    .io_1(Delay_Pipe_Hw_3_io_1),
    .io_0(Delay_Pipe_Hw_3_io_0)
  );
  Delay_Pipe_Hw_1 Delay_Pipe_Hw_4 ( // @[Dedicated_PE.scala 86:39:@4234.4]
    .clock(Delay_Pipe_Hw_4_clock),
    .reset(Delay_Pipe_Hw_4_reset),
    .io_2(Delay_Pipe_Hw_4_io_2),
    .io_1(Delay_Pipe_Hw_4_io_1),
    .io_0(Delay_Pipe_Hw_4_io_0)
  );
  Delay_Pipe_Hw_1 Delay_Pipe_Hw_5 ( // @[Dedicated_PE.scala 86:39:@4237.4]
    .clock(Delay_Pipe_Hw_5_clock),
    .reset(Delay_Pipe_Hw_5_reset),
    .io_2(Delay_Pipe_Hw_5_io_2),
    .io_1(Delay_Pipe_Hw_5_io_1),
    .io_0(Delay_Pipe_Hw_5_io_0)
  );
  Arithmetic_Logic_Unit_Hw Arithmetic_Logic_Unit_Hw_1 ( // @[Dedicated_PE.scala 85:32:@4240.4]
    .clock(Arithmetic_Logic_Unit_Hw_1_clock),
    .reset(Arithmetic_Logic_Unit_Hw_1_reset),
    .io_4(Arithmetic_Logic_Unit_Hw_1_io_4),
    .io_3(Arithmetic_Logic_Unit_Hw_1_io_3),
    .io_2(Arithmetic_Logic_Unit_Hw_1_io_2),
    .io_1(Arithmetic_Logic_Unit_Hw_1_io_1),
    .io_0(Arithmetic_Logic_Unit_Hw_1_io_0)
  );
  Delay_Pipe_Hw_6 Delay_Pipe_Hw_6 ( // @[Dedicated_PE.scala 86:39:@4243.4]
    .clock(Delay_Pipe_Hw_6_clock),
    .reset(Delay_Pipe_Hw_6_reset),
    .io_2(Delay_Pipe_Hw_6_io_2),
    .io_1(Delay_Pipe_Hw_6_io_1),
    .io_0(Delay_Pipe_Hw_6_io_0)
  );
  Delay_Pipe_Hw_7 Delay_Pipe_Hw_7 ( // @[Dedicated_PE.scala 86:39:@4246.4]
    .clock(Delay_Pipe_Hw_7_clock),
    .reset(Delay_Pipe_Hw_7_reset),
    .io_2(Delay_Pipe_Hw_7_io_2),
    .io_1(Delay_Pipe_Hw_7_io_1),
    .io_0(Delay_Pipe_Hw_7_io_0)
  );
  Delay_Pipe_Hw_7 Delay_Pipe_Hw_8 ( // @[Dedicated_PE.scala 86:39:@4249.4]
    .clock(Delay_Pipe_Hw_8_clock),
    .reset(Delay_Pipe_Hw_8_reset),
    .io_2(Delay_Pipe_Hw_8_io_2),
    .io_1(Delay_Pipe_Hw_8_io_1),
    .io_0(Delay_Pipe_Hw_8_io_0)
  );
  Arithmetic_Logic_Unit_Hw_2 Arithmetic_Logic_Unit_Hw_2 ( // @[Dedicated_PE.scala 85:32:@4252.4]
    .clock(Arithmetic_Logic_Unit_Hw_2_clock),
    .reset(Arithmetic_Logic_Unit_Hw_2_reset),
    .io_4(Arithmetic_Logic_Unit_Hw_2_io_4),
    .io_3(Arithmetic_Logic_Unit_Hw_2_io_3),
    .io_2(Arithmetic_Logic_Unit_Hw_2_io_2),
    .io_1(Arithmetic_Logic_Unit_Hw_2_io_1),
    .io_0(Arithmetic_Logic_Unit_Hw_2_io_0)
  );
  Delay_Pipe_Hw_6 Delay_Pipe_Hw_9 ( // @[Dedicated_PE.scala 86:39:@4255.4]
    .clock(Delay_Pipe_Hw_9_clock),
    .reset(Delay_Pipe_Hw_9_reset),
    .io_2(Delay_Pipe_Hw_9_io_2),
    .io_1(Delay_Pipe_Hw_9_io_1),
    .io_0(Delay_Pipe_Hw_9_io_0)
  );
  Delay_Pipe_Hw_7 Delay_Pipe_Hw_10 ( // @[Dedicated_PE.scala 86:39:@4258.4]
    .clock(Delay_Pipe_Hw_10_clock),
    .reset(Delay_Pipe_Hw_10_reset),
    .io_2(Delay_Pipe_Hw_10_io_2),
    .io_1(Delay_Pipe_Hw_10_io_1),
    .io_0(Delay_Pipe_Hw_10_io_0)
  );
  Delay_Pipe_Hw_7 Delay_Pipe_Hw_11 ( // @[Dedicated_PE.scala 86:39:@4261.4]
    .clock(Delay_Pipe_Hw_11_clock),
    .reset(Delay_Pipe_Hw_11_reset),
    .io_2(Delay_Pipe_Hw_11_io_2),
    .io_1(Delay_Pipe_Hw_11_io_1),
    .io_0(Delay_Pipe_Hw_11_io_0)
  );
  Arithmetic_Logic_Unit_Hw_2 Arithmetic_Logic_Unit_Hw_3 ( // @[Dedicated_PE.scala 85:32:@4264.4]
    .clock(Arithmetic_Logic_Unit_Hw_3_clock),
    .reset(Arithmetic_Logic_Unit_Hw_3_reset),
    .io_4(Arithmetic_Logic_Unit_Hw_3_io_4),
    .io_3(Arithmetic_Logic_Unit_Hw_3_io_3),
    .io_2(Arithmetic_Logic_Unit_Hw_3_io_2),
    .io_1(Arithmetic_Logic_Unit_Hw_3_io_1),
    .io_0(Arithmetic_Logic_Unit_Hw_3_io_0)
  );
  Delay_Pipe_Hw_6 Delay_Pipe_Hw_12 ( // @[Dedicated_PE.scala 86:39:@4267.4]
    .clock(Delay_Pipe_Hw_12_clock),
    .reset(Delay_Pipe_Hw_12_reset),
    .io_2(Delay_Pipe_Hw_12_io_2),
    .io_1(Delay_Pipe_Hw_12_io_1),
    .io_0(Delay_Pipe_Hw_12_io_0)
  );
  Delay_Pipe_Hw_7 Delay_Pipe_Hw_13 ( // @[Dedicated_PE.scala 86:39:@4270.4]
    .clock(Delay_Pipe_Hw_13_clock),
    .reset(Delay_Pipe_Hw_13_reset),
    .io_2(Delay_Pipe_Hw_13_io_2),
    .io_1(Delay_Pipe_Hw_13_io_1),
    .io_0(Delay_Pipe_Hw_13_io_0)
  );
  Delay_Pipe_Hw_7 Delay_Pipe_Hw_14 ( // @[Dedicated_PE.scala 86:39:@4273.4]
    .clock(Delay_Pipe_Hw_14_clock),
    .reset(Delay_Pipe_Hw_14_reset),
    .io_2(Delay_Pipe_Hw_14_io_2),
    .io_1(Delay_Pipe_Hw_14_io_1),
    .io_0(Delay_Pipe_Hw_14_io_0)
  );
  Arithmetic_Logic_Unit_Hw_2 Arithmetic_Logic_Unit_Hw_4 ( // @[Dedicated_PE.scala 85:32:@4276.4]
    .clock(Arithmetic_Logic_Unit_Hw_4_clock),
    .reset(Arithmetic_Logic_Unit_Hw_4_reset),
    .io_4(Arithmetic_Logic_Unit_Hw_4_io_4),
    .io_3(Arithmetic_Logic_Unit_Hw_4_io_3),
    .io_2(Arithmetic_Logic_Unit_Hw_4_io_2),
    .io_1(Arithmetic_Logic_Unit_Hw_4_io_1),
    .io_0(Arithmetic_Logic_Unit_Hw_4_io_0)
  );
  Delay_Pipe_Hw_6 Delay_Pipe_Hw_15 ( // @[Dedicated_PE.scala 86:39:@4279.4]
    .clock(Delay_Pipe_Hw_15_clock),
    .reset(Delay_Pipe_Hw_15_reset),
    .io_2(Delay_Pipe_Hw_15_io_2),
    .io_1(Delay_Pipe_Hw_15_io_1),
    .io_0(Delay_Pipe_Hw_15_io_0)
  );
  Delay_Pipe_Hw_7 Delay_Pipe_Hw_16 ( // @[Dedicated_PE.scala 86:39:@4282.4]
    .clock(Delay_Pipe_Hw_16_clock),
    .reset(Delay_Pipe_Hw_16_reset),
    .io_2(Delay_Pipe_Hw_16_io_2),
    .io_1(Delay_Pipe_Hw_16_io_1),
    .io_0(Delay_Pipe_Hw_16_io_0)
  );
  Delay_Pipe_Hw_7 Delay_Pipe_Hw_17 ( // @[Dedicated_PE.scala 86:39:@4285.4]
    .clock(Delay_Pipe_Hw_17_clock),
    .reset(Delay_Pipe_Hw_17_reset),
    .io_2(Delay_Pipe_Hw_17_io_2),
    .io_1(Delay_Pipe_Hw_17_io_1),
    .io_0(Delay_Pipe_Hw_17_io_0)
  );
  Arithmetic_Logic_Unit_Hw_2 Arithmetic_Logic_Unit_Hw_5 ( // @[Dedicated_PE.scala 85:32:@4288.4]
    .clock(Arithmetic_Logic_Unit_Hw_5_clock),
    .reset(Arithmetic_Logic_Unit_Hw_5_reset),
    .io_4(Arithmetic_Logic_Unit_Hw_5_io_4),
    .io_3(Arithmetic_Logic_Unit_Hw_5_io_3),
    .io_2(Arithmetic_Logic_Unit_Hw_5_io_2),
    .io_1(Arithmetic_Logic_Unit_Hw_5_io_1),
    .io_0(Arithmetic_Logic_Unit_Hw_5_io_0)
  );
  Multiplexer_Hw Multiplexer_Hw ( // @[Dedicated_PE.scala 84:32:@4291.4]
    .io_4(Multiplexer_Hw_io_4),
    .io_3(Multiplexer_Hw_io_3),
    .io_2(Multiplexer_Hw_io_2),
    .io_1(Multiplexer_Hw_io_1),
    .io_0(Multiplexer_Hw_io_0)
  );
  Multiplexer_Hw Multiplexer_Hw_1 ( // @[Dedicated_PE.scala 84:32:@4294.4]
    .io_4(Multiplexer_Hw_1_io_4),
    .io_3(Multiplexer_Hw_1_io_3),
    .io_2(Multiplexer_Hw_1_io_2),
    .io_1(Multiplexer_Hw_1_io_1),
    .io_0(Multiplexer_Hw_1_io_0)
  );
  Multiplexer_Hw Multiplexer_Hw_2 ( // @[Dedicated_PE.scala 84:32:@4297.4]
    .io_4(Multiplexer_Hw_2_io_4),
    .io_3(Multiplexer_Hw_2_io_3),
    .io_2(Multiplexer_Hw_2_io_2),
    .io_1(Multiplexer_Hw_2_io_1),
    .io_0(Multiplexer_Hw_2_io_0)
  );
  Multiplexer_Hw Multiplexer_Hw_3 ( // @[Dedicated_PE.scala 84:32:@4300.4]
    .io_4(Multiplexer_Hw_3_io_4),
    .io_3(Multiplexer_Hw_3_io_3),
    .io_2(Multiplexer_Hw_3_io_2),
    .io_1(Multiplexer_Hw_3_io_1),
    .io_0(Multiplexer_Hw_3_io_0)
  );
  Multiplexer_Hw Multiplexer_Hw_4 ( // @[Dedicated_PE.scala 84:32:@4303.4]
    .io_4(Multiplexer_Hw_4_io_4),
    .io_3(Multiplexer_Hw_4_io_3),
    .io_2(Multiplexer_Hw_4_io_2),
    .io_1(Multiplexer_Hw_4_io_1),
    .io_0(Multiplexer_Hw_4_io_0)
  );
  Multiplexer_Hw Multiplexer_Hw_5 ( // @[Dedicated_PE.scala 84:32:@4306.4]
    .io_4(Multiplexer_Hw_5_io_4),
    .io_3(Multiplexer_Hw_5_io_3),
    .io_2(Multiplexer_Hw_5_io_2),
    .io_1(Multiplexer_Hw_5_io_1),
    .io_0(Multiplexer_Hw_5_io_0)
  );
  Multiplexer_Hw_6 Multiplexer_Hw_6 ( // @[Dedicated_PE.scala 84:32:@4309.4]
    .io_4(Multiplexer_Hw_6_io_4),
    .io_3(Multiplexer_Hw_6_io_3),
    .io_2(Multiplexer_Hw_6_io_2),
    .io_1(Multiplexer_Hw_6_io_1),
    .io_0(Multiplexer_Hw_6_io_0)
  );
  Multiplexer_Hw_6 Multiplexer_Hw_7 ( // @[Dedicated_PE.scala 84:32:@4312.4]
    .io_4(Multiplexer_Hw_7_io_4),
    .io_3(Multiplexer_Hw_7_io_3),
    .io_2(Multiplexer_Hw_7_io_2),
    .io_1(Multiplexer_Hw_7_io_1),
    .io_0(Multiplexer_Hw_7_io_0)
  );
  Multiplexer_Hw_6 Multiplexer_Hw_8 ( // @[Dedicated_PE.scala 84:32:@4315.4]
    .io_4(Multiplexer_Hw_8_io_4),
    .io_3(Multiplexer_Hw_8_io_3),
    .io_2(Multiplexer_Hw_8_io_2),
    .io_1(Multiplexer_Hw_8_io_1),
    .io_0(Multiplexer_Hw_8_io_0)
  );
  Multiplexer_Hw_6 Multiplexer_Hw_9 ( // @[Dedicated_PE.scala 84:32:@4318.4]
    .io_4(Multiplexer_Hw_9_io_4),
    .io_3(Multiplexer_Hw_9_io_3),
    .io_2(Multiplexer_Hw_9_io_2),
    .io_1(Multiplexer_Hw_9_io_1),
    .io_0(Multiplexer_Hw_9_io_0)
  );
  Multiplexer_Hw_6 Multiplexer_Hw_10 ( // @[Dedicated_PE.scala 84:32:@4321.4]
    .io_4(Multiplexer_Hw_10_io_4),
    .io_3(Multiplexer_Hw_10_io_3),
    .io_2(Multiplexer_Hw_10_io_2),
    .io_1(Multiplexer_Hw_10_io_1),
    .io_0(Multiplexer_Hw_10_io_0)
  );
  Multiplexer_Hw_6 Multiplexer_Hw_11 ( // @[Dedicated_PE.scala 84:32:@4324.4]
    .io_4(Multiplexer_Hw_11_io_4),
    .io_3(Multiplexer_Hw_11_io_3),
    .io_2(Multiplexer_Hw_11_io_2),
    .io_1(Multiplexer_Hw_11_io_1),
    .io_0(Multiplexer_Hw_11_io_0)
  );
  Multiplexer_Hw_6 Multiplexer_Hw_12 ( // @[Dedicated_PE.scala 84:32:@4327.4]
    .io_4(Multiplexer_Hw_12_io_4),
    .io_3(Multiplexer_Hw_12_io_3),
    .io_2(Multiplexer_Hw_12_io_2),
    .io_1(Multiplexer_Hw_12_io_1),
    .io_0(Multiplexer_Hw_12_io_0)
  );
  Multiplexer_Hw_6 Multiplexer_Hw_13 ( // @[Dedicated_PE.scala 84:32:@4330.4]
    .io_4(Multiplexer_Hw_13_io_4),
    .io_3(Multiplexer_Hw_13_io_3),
    .io_2(Multiplexer_Hw_13_io_2),
    .io_1(Multiplexer_Hw_13_io_1),
    .io_0(Multiplexer_Hw_13_io_0)
  );
  Multiplexer_Hw_6 Multiplexer_Hw_14 ( // @[Dedicated_PE.scala 84:32:@4333.4]
    .io_4(Multiplexer_Hw_14_io_4),
    .io_3(Multiplexer_Hw_14_io_3),
    .io_2(Multiplexer_Hw_14_io_2),
    .io_1(Multiplexer_Hw_14_io_1),
    .io_0(Multiplexer_Hw_14_io_0)
  );
  Multiplexer_Hw_6 Multiplexer_Hw_15 ( // @[Dedicated_PE.scala 84:32:@4336.4]
    .io_4(Multiplexer_Hw_15_io_4),
    .io_3(Multiplexer_Hw_15_io_3),
    .io_2(Multiplexer_Hw_15_io_2),
    .io_1(Multiplexer_Hw_15_io_1),
    .io_0(Multiplexer_Hw_15_io_0)
  );
  Multiplexer_Hw_6 Multiplexer_Hw_16 ( // @[Dedicated_PE.scala 84:32:@4339.4]
    .io_4(Multiplexer_Hw_16_io_4),
    .io_3(Multiplexer_Hw_16_io_3),
    .io_2(Multiplexer_Hw_16_io_2),
    .io_1(Multiplexer_Hw_16_io_1),
    .io_0(Multiplexer_Hw_16_io_0)
  );
  Multiplexer_Hw_6 Multiplexer_Hw_17 ( // @[Dedicated_PE.scala 84:32:@4342.4]
    .io_4(Multiplexer_Hw_17_io_4),
    .io_3(Multiplexer_Hw_17_io_3),
    .io_2(Multiplexer_Hw_17_io_2),
    .io_1(Multiplexer_Hw_17_io_1),
    .io_0(Multiplexer_Hw_17_io_0)
  );
  assign _T_167 = io_24_write_index[2:0]; // @[:@4526.6]
  assign _GEN_0 = 3'h0 == _T_167 ? io_24_write_data : config_registers_0; // @[Dedicated_PE.scala 137:47:@4527.6]
  assign _GEN_1 = 3'h1 == _T_167 ? io_24_write_data : config_registers_1; // @[Dedicated_PE.scala 137:47:@4527.6]
  assign _GEN_2 = 3'h2 == _T_167 ? io_24_write_data : config_registers_2; // @[Dedicated_PE.scala 137:47:@4527.6]
  assign _GEN_3 = 3'h3 == _T_167 ? io_24_write_data : config_registers_3; // @[Dedicated_PE.scala 137:47:@4527.6]
  assign _GEN_4 = 3'h4 == _T_167 ? io_24_write_data : config_registers_4; // @[Dedicated_PE.scala 137:47:@4527.6]
  assign _GEN_5 = 3'h5 == _T_167 ? io_24_write_data : config_registers_5; // @[Dedicated_PE.scala 137:47:@4527.6]
  assign _GEN_6 = 3'h6 == _T_167 ? io_24_write_data : config_registers_6; // @[Dedicated_PE.scala 137:47:@4527.6]
  assign _GEN_7 = 3'h7 == _T_167 ? io_24_write_data : config_registers_7; // @[Dedicated_PE.scala 137:47:@4527.6]
  assign io_24_read_ack = 1'h0; // @[Dedicated_PE.scala 140:24:@4530.4]
  assign io_24_read_data = 16'h0; // @[Dedicated_PE.scala 141:25:@4531.4]
  assign io_24_write_ack = 1'h1; // @[Dedicated_PE.scala 139:25:@4529.4]
  assign io_23 = Arithmetic_Logic_Unit_Hw_5_io_2; // @[Dedicated_PE.scala 121:15:@4368.4]
  assign io_22 = Arithmetic_Logic_Unit_Hw_4_io_2; // @[Dedicated_PE.scala 121:15:@4364.4]
  assign io_21 = Arithmetic_Logic_Unit_Hw_3_io_2; // @[Dedicated_PE.scala 121:15:@4360.4]
  assign io_20 = Arithmetic_Logic_Unit_Hw_2_io_2; // @[Dedicated_PE.scala 121:15:@4356.4]
  assign io_19 = Arithmetic_Logic_Unit_Hw_1_io_2; // @[Dedicated_PE.scala 121:15:@4352.4]
  assign io_18 = Arithmetic_Logic_Unit_Hw_io_2; // @[Dedicated_PE.scala 121:15:@4348.4]
  assign Delay_Pipe_Hw_clock = clock; // @[:@4220.4]
  assign Delay_Pipe_Hw_reset = reset; // @[:@4221.4]
  assign Delay_Pipe_Hw_io_2 = config_registers_0[2:0]; // @[Dedicated_PE.scala 130:45:@4442.4]
  assign Delay_Pipe_Hw_io_0 = Multiplexer_Hw_io_3; // @[Dedicated_PE.scala 121:15:@4372.4]
  assign Delay_Pipe_Hw_1_clock = clock; // @[:@4223.4]
  assign Delay_Pipe_Hw_1_reset = reset; // @[:@4224.4]
  assign Delay_Pipe_Hw_1_io_2 = config_registers_0[4:3]; // @[Dedicated_PE.scala 130:45:@4444.4]
  assign Delay_Pipe_Hw_1_io_0 = Multiplexer_Hw_1_io_3; // @[Dedicated_PE.scala 121:15:@4376.4]
  assign Delay_Pipe_Hw_2_clock = clock; // @[:@4226.4]
  assign Delay_Pipe_Hw_2_reset = reset; // @[:@4227.4]
  assign Delay_Pipe_Hw_2_io_2 = config_registers_0[6:5]; // @[Dedicated_PE.scala 130:45:@4446.4]
  assign Delay_Pipe_Hw_2_io_0 = Multiplexer_Hw_2_io_3; // @[Dedicated_PE.scala 121:15:@4380.4]
  assign Arithmetic_Logic_Unit_Hw_clock = clock; // @[:@4229.4]
  assign Arithmetic_Logic_Unit_Hw_reset = reset; // @[:@4230.4]
  assign Arithmetic_Logic_Unit_Hw_io_4 = config_registers_0[11:7]; // @[Dedicated_PE.scala 130:45:@4448.4]
  assign Arithmetic_Logic_Unit_Hw_io_3 = Delay_Pipe_Hw_2_io_1; // @[Dedicated_PE.scala 121:15:@4347.4]
  assign Arithmetic_Logic_Unit_Hw_io_1 = Delay_Pipe_Hw_1_io_1; // @[Dedicated_PE.scala 121:15:@4346.4]
  assign Arithmetic_Logic_Unit_Hw_io_0 = Delay_Pipe_Hw_io_1; // @[Dedicated_PE.scala 121:15:@4345.4]
  assign Delay_Pipe_Hw_3_clock = clock; // @[:@4232.4]
  assign Delay_Pipe_Hw_3_reset = reset; // @[:@4233.4]
  assign Delay_Pipe_Hw_3_io_2 = config_registers_0[14:12]; // @[Dedicated_PE.scala 130:45:@4450.4]
  assign Delay_Pipe_Hw_3_io_0 = Multiplexer_Hw_3_io_3; // @[Dedicated_PE.scala 121:15:@4384.4]
  assign Delay_Pipe_Hw_4_clock = clock; // @[:@4235.4]
  assign Delay_Pipe_Hw_4_reset = reset; // @[:@4236.4]
  assign Delay_Pipe_Hw_4_io_2 = config_registers_1[1:0]; // @[Dedicated_PE.scala 130:45:@4452.4]
  assign Delay_Pipe_Hw_4_io_0 = Multiplexer_Hw_4_io_3; // @[Dedicated_PE.scala 121:15:@4388.4]
  assign Delay_Pipe_Hw_5_clock = clock; // @[:@4238.4]
  assign Delay_Pipe_Hw_5_reset = reset; // @[:@4239.4]
  assign Delay_Pipe_Hw_5_io_2 = config_registers_1[3:2]; // @[Dedicated_PE.scala 130:45:@4454.4]
  assign Delay_Pipe_Hw_5_io_0 = Multiplexer_Hw_5_io_3; // @[Dedicated_PE.scala 121:15:@4392.4]
  assign Arithmetic_Logic_Unit_Hw_1_clock = clock; // @[:@4241.4]
  assign Arithmetic_Logic_Unit_Hw_1_reset = reset; // @[:@4242.4]
  assign Arithmetic_Logic_Unit_Hw_1_io_4 = config_registers_1[8:4]; // @[Dedicated_PE.scala 130:45:@4456.4]
  assign Arithmetic_Logic_Unit_Hw_1_io_3 = Delay_Pipe_Hw_5_io_1; // @[Dedicated_PE.scala 121:15:@4351.4]
  assign Arithmetic_Logic_Unit_Hw_1_io_1 = Delay_Pipe_Hw_4_io_1; // @[Dedicated_PE.scala 121:15:@4350.4]
  assign Arithmetic_Logic_Unit_Hw_1_io_0 = Delay_Pipe_Hw_3_io_1; // @[Dedicated_PE.scala 121:15:@4349.4]
  assign Delay_Pipe_Hw_6_clock = clock; // @[:@4244.4]
  assign Delay_Pipe_Hw_6_reset = reset; // @[:@4245.4]
  assign Delay_Pipe_Hw_6_io_2 = config_registers_1[11:9]; // @[Dedicated_PE.scala 130:45:@4458.4]
  assign Delay_Pipe_Hw_6_io_0 = Multiplexer_Hw_6_io_3; // @[Dedicated_PE.scala 121:15:@4396.4]
  assign Delay_Pipe_Hw_7_clock = clock; // @[:@4247.4]
  assign Delay_Pipe_Hw_7_reset = reset; // @[:@4248.4]
  assign Delay_Pipe_Hw_7_io_2 = config_registers_1[13:12]; // @[Dedicated_PE.scala 130:45:@4460.4]
  assign Delay_Pipe_Hw_7_io_0 = Multiplexer_Hw_7_io_3; // @[Dedicated_PE.scala 121:15:@4400.4]
  assign Delay_Pipe_Hw_8_clock = clock; // @[:@4250.4]
  assign Delay_Pipe_Hw_8_reset = reset; // @[:@4251.4]
  assign Delay_Pipe_Hw_8_io_2 = config_registers_1[15:14]; // @[Dedicated_PE.scala 130:45:@4462.4]
  assign Delay_Pipe_Hw_8_io_0 = Multiplexer_Hw_8_io_3; // @[Dedicated_PE.scala 121:15:@4404.4]
  assign Arithmetic_Logic_Unit_Hw_2_clock = clock; // @[:@4253.4]
  assign Arithmetic_Logic_Unit_Hw_2_reset = reset; // @[:@4254.4]
  assign Arithmetic_Logic_Unit_Hw_2_io_4 = config_registers_2[4:0]; // @[Dedicated_PE.scala 130:45:@4464.4]
  assign Arithmetic_Logic_Unit_Hw_2_io_3 = Delay_Pipe_Hw_8_io_1; // @[Dedicated_PE.scala 121:15:@4355.4]
  assign Arithmetic_Logic_Unit_Hw_2_io_1 = Delay_Pipe_Hw_7_io_1; // @[Dedicated_PE.scala 121:15:@4354.4]
  assign Arithmetic_Logic_Unit_Hw_2_io_0 = Delay_Pipe_Hw_6_io_1; // @[Dedicated_PE.scala 121:15:@4353.4]
  assign Delay_Pipe_Hw_9_clock = clock; // @[:@4256.4]
  assign Delay_Pipe_Hw_9_reset = reset; // @[:@4257.4]
  assign Delay_Pipe_Hw_9_io_2 = config_registers_2[7:5]; // @[Dedicated_PE.scala 130:45:@4466.4]
  assign Delay_Pipe_Hw_9_io_0 = Multiplexer_Hw_9_io_3; // @[Dedicated_PE.scala 121:15:@4408.4]
  assign Delay_Pipe_Hw_10_clock = clock; // @[:@4259.4]
  assign Delay_Pipe_Hw_10_reset = reset; // @[:@4260.4]
  assign Delay_Pipe_Hw_10_io_2 = config_registers_2[9:8]; // @[Dedicated_PE.scala 130:45:@4468.4]
  assign Delay_Pipe_Hw_10_io_0 = Multiplexer_Hw_10_io_3; // @[Dedicated_PE.scala 121:15:@4412.4]
  assign Delay_Pipe_Hw_11_clock = clock; // @[:@4262.4]
  assign Delay_Pipe_Hw_11_reset = reset; // @[:@4263.4]
  assign Delay_Pipe_Hw_11_io_2 = config_registers_2[11:10]; // @[Dedicated_PE.scala 130:45:@4470.4]
  assign Delay_Pipe_Hw_11_io_0 = Multiplexer_Hw_11_io_3; // @[Dedicated_PE.scala 121:15:@4416.4]
  assign Arithmetic_Logic_Unit_Hw_3_clock = clock; // @[:@4265.4]
  assign Arithmetic_Logic_Unit_Hw_3_reset = reset; // @[:@4266.4]
  assign Arithmetic_Logic_Unit_Hw_3_io_4 = config_registers_3[4:0]; // @[Dedicated_PE.scala 130:45:@4472.4]
  assign Arithmetic_Logic_Unit_Hw_3_io_3 = Delay_Pipe_Hw_11_io_1; // @[Dedicated_PE.scala 121:15:@4359.4]
  assign Arithmetic_Logic_Unit_Hw_3_io_1 = Delay_Pipe_Hw_10_io_1; // @[Dedicated_PE.scala 121:15:@4358.4]
  assign Arithmetic_Logic_Unit_Hw_3_io_0 = Delay_Pipe_Hw_9_io_1; // @[Dedicated_PE.scala 121:15:@4357.4]
  assign Delay_Pipe_Hw_12_clock = clock; // @[:@4268.4]
  assign Delay_Pipe_Hw_12_reset = reset; // @[:@4269.4]
  assign Delay_Pipe_Hw_12_io_2 = config_registers_3[7:5]; // @[Dedicated_PE.scala 130:45:@4474.4]
  assign Delay_Pipe_Hw_12_io_0 = Multiplexer_Hw_12_io_3; // @[Dedicated_PE.scala 121:15:@4420.4]
  assign Delay_Pipe_Hw_13_clock = clock; // @[:@4271.4]
  assign Delay_Pipe_Hw_13_reset = reset; // @[:@4272.4]
  assign Delay_Pipe_Hw_13_io_2 = config_registers_3[9:8]; // @[Dedicated_PE.scala 130:45:@4476.4]
  assign Delay_Pipe_Hw_13_io_0 = Multiplexer_Hw_13_io_3; // @[Dedicated_PE.scala 121:15:@4424.4]
  assign Delay_Pipe_Hw_14_clock = clock; // @[:@4274.4]
  assign Delay_Pipe_Hw_14_reset = reset; // @[:@4275.4]
  assign Delay_Pipe_Hw_14_io_2 = config_registers_3[11:10]; // @[Dedicated_PE.scala 130:45:@4478.4]
  assign Delay_Pipe_Hw_14_io_0 = Multiplexer_Hw_14_io_3; // @[Dedicated_PE.scala 121:15:@4428.4]
  assign Arithmetic_Logic_Unit_Hw_4_clock = clock; // @[:@4277.4]
  assign Arithmetic_Logic_Unit_Hw_4_reset = reset; // @[:@4278.4]
  assign Arithmetic_Logic_Unit_Hw_4_io_4 = config_registers_4[4:0]; // @[Dedicated_PE.scala 130:45:@4480.4]
  assign Arithmetic_Logic_Unit_Hw_4_io_3 = Delay_Pipe_Hw_14_io_1; // @[Dedicated_PE.scala 121:15:@4363.4]
  assign Arithmetic_Logic_Unit_Hw_4_io_1 = Delay_Pipe_Hw_13_io_1; // @[Dedicated_PE.scala 121:15:@4362.4]
  assign Arithmetic_Logic_Unit_Hw_4_io_0 = Delay_Pipe_Hw_12_io_1; // @[Dedicated_PE.scala 121:15:@4361.4]
  assign Delay_Pipe_Hw_15_clock = clock; // @[:@4280.4]
  assign Delay_Pipe_Hw_15_reset = reset; // @[:@4281.4]
  assign Delay_Pipe_Hw_15_io_2 = config_registers_4[7:5]; // @[Dedicated_PE.scala 130:45:@4482.4]
  assign Delay_Pipe_Hw_15_io_0 = Multiplexer_Hw_15_io_3; // @[Dedicated_PE.scala 121:15:@4432.4]
  assign Delay_Pipe_Hw_16_clock = clock; // @[:@4283.4]
  assign Delay_Pipe_Hw_16_reset = reset; // @[:@4284.4]
  assign Delay_Pipe_Hw_16_io_2 = config_registers_4[9:8]; // @[Dedicated_PE.scala 130:45:@4484.4]
  assign Delay_Pipe_Hw_16_io_0 = Multiplexer_Hw_16_io_3; // @[Dedicated_PE.scala 121:15:@4436.4]
  assign Delay_Pipe_Hw_17_clock = clock; // @[:@4286.4]
  assign Delay_Pipe_Hw_17_reset = reset; // @[:@4287.4]
  assign Delay_Pipe_Hw_17_io_2 = config_registers_4[11:10]; // @[Dedicated_PE.scala 130:45:@4486.4]
  assign Delay_Pipe_Hw_17_io_0 = Multiplexer_Hw_17_io_3; // @[Dedicated_PE.scala 121:15:@4440.4]
  assign Arithmetic_Logic_Unit_Hw_5_clock = clock; // @[:@4289.4]
  assign Arithmetic_Logic_Unit_Hw_5_reset = reset; // @[:@4290.4]
  assign Arithmetic_Logic_Unit_Hw_5_io_4 = config_registers_5[4:0]; // @[Dedicated_PE.scala 130:45:@4488.4]
  assign Arithmetic_Logic_Unit_Hw_5_io_3 = Delay_Pipe_Hw_17_io_1; // @[Dedicated_PE.scala 121:15:@4367.4]
  assign Arithmetic_Logic_Unit_Hw_5_io_1 = Delay_Pipe_Hw_16_io_1; // @[Dedicated_PE.scala 121:15:@4366.4]
  assign Arithmetic_Logic_Unit_Hw_5_io_0 = Delay_Pipe_Hw_15_io_1; // @[Dedicated_PE.scala 121:15:@4365.4]
  assign Multiplexer_Hw_io_4 = config_registers_5[6:5]; // @[Dedicated_PE.scala 130:45:@4490.4]
  assign Multiplexer_Hw_io_2 = io_4; // @[Dedicated_PE.scala 121:15:@4371.4]
  assign Multiplexer_Hw_io_1 = io_2; // @[Dedicated_PE.scala 121:15:@4370.4]
  assign Multiplexer_Hw_io_0 = io_0; // @[Dedicated_PE.scala 121:15:@4369.4]
  assign Multiplexer_Hw_1_io_4 = config_registers_5[8:7]; // @[Dedicated_PE.scala 130:45:@4492.4]
  assign Multiplexer_Hw_1_io_2 = io_4; // @[Dedicated_PE.scala 121:15:@4375.4]
  assign Multiplexer_Hw_1_io_1 = io_2; // @[Dedicated_PE.scala 121:15:@4374.4]
  assign Multiplexer_Hw_1_io_0 = io_0; // @[Dedicated_PE.scala 121:15:@4373.4]
  assign Multiplexer_Hw_2_io_4 = config_registers_5[10:9]; // @[Dedicated_PE.scala 130:45:@4494.4]
  assign Multiplexer_Hw_2_io_2 = io_4; // @[Dedicated_PE.scala 121:15:@4379.4]
  assign Multiplexer_Hw_2_io_1 = io_2; // @[Dedicated_PE.scala 121:15:@4378.4]
  assign Multiplexer_Hw_2_io_0 = io_0; // @[Dedicated_PE.scala 121:15:@4377.4]
  assign Multiplexer_Hw_3_io_4 = config_registers_5[12:11]; // @[Dedicated_PE.scala 130:45:@4496.4]
  assign Multiplexer_Hw_3_io_2 = io_5; // @[Dedicated_PE.scala 121:15:@4383.4]
  assign Multiplexer_Hw_3_io_1 = io_3; // @[Dedicated_PE.scala 121:15:@4382.4]
  assign Multiplexer_Hw_3_io_0 = io_1; // @[Dedicated_PE.scala 121:15:@4381.4]
  assign Multiplexer_Hw_4_io_4 = config_registers_5[14:13]; // @[Dedicated_PE.scala 130:45:@4498.4]
  assign Multiplexer_Hw_4_io_2 = io_5; // @[Dedicated_PE.scala 121:15:@4387.4]
  assign Multiplexer_Hw_4_io_1 = io_3; // @[Dedicated_PE.scala 121:15:@4386.4]
  assign Multiplexer_Hw_4_io_0 = io_1; // @[Dedicated_PE.scala 121:15:@4385.4]
  assign Multiplexer_Hw_5_io_4 = config_registers_6[1:0]; // @[Dedicated_PE.scala 130:45:@4500.4]
  assign Multiplexer_Hw_5_io_2 = io_5; // @[Dedicated_PE.scala 121:15:@4391.4]
  assign Multiplexer_Hw_5_io_1 = io_3; // @[Dedicated_PE.scala 121:15:@4390.4]
  assign Multiplexer_Hw_5_io_0 = io_1; // @[Dedicated_PE.scala 121:15:@4389.4]
  assign Multiplexer_Hw_6_io_4 = config_registers_6[3:2]; // @[Dedicated_PE.scala 130:45:@4502.4]
  assign Multiplexer_Hw_6_io_2 = io_14; // @[Dedicated_PE.scala 121:15:@4395.4]
  assign Multiplexer_Hw_6_io_1 = io_10; // @[Dedicated_PE.scala 121:15:@4394.4]
  assign Multiplexer_Hw_6_io_0 = io_6; // @[Dedicated_PE.scala 121:15:@4393.4]
  assign Multiplexer_Hw_7_io_4 = config_registers_6[5:4]; // @[Dedicated_PE.scala 130:45:@4504.4]
  assign Multiplexer_Hw_7_io_2 = io_14; // @[Dedicated_PE.scala 121:15:@4399.4]
  assign Multiplexer_Hw_7_io_1 = io_10; // @[Dedicated_PE.scala 121:15:@4398.4]
  assign Multiplexer_Hw_7_io_0 = io_6; // @[Dedicated_PE.scala 121:15:@4397.4]
  assign Multiplexer_Hw_8_io_4 = config_registers_6[7:6]; // @[Dedicated_PE.scala 130:45:@4506.4]
  assign Multiplexer_Hw_8_io_2 = io_14; // @[Dedicated_PE.scala 121:15:@4403.4]
  assign Multiplexer_Hw_8_io_1 = io_10; // @[Dedicated_PE.scala 121:15:@4402.4]
  assign Multiplexer_Hw_8_io_0 = io_6; // @[Dedicated_PE.scala 121:15:@4401.4]
  assign Multiplexer_Hw_9_io_4 = config_registers_6[9:8]; // @[Dedicated_PE.scala 130:45:@4508.4]
  assign Multiplexer_Hw_9_io_2 = io_15; // @[Dedicated_PE.scala 121:15:@4407.4]
  assign Multiplexer_Hw_9_io_1 = io_11; // @[Dedicated_PE.scala 121:15:@4406.4]
  assign Multiplexer_Hw_9_io_0 = io_7; // @[Dedicated_PE.scala 121:15:@4405.4]
  assign Multiplexer_Hw_10_io_4 = config_registers_6[11:10]; // @[Dedicated_PE.scala 130:45:@4510.4]
  assign Multiplexer_Hw_10_io_2 = io_15; // @[Dedicated_PE.scala 121:15:@4411.4]
  assign Multiplexer_Hw_10_io_1 = io_11; // @[Dedicated_PE.scala 121:15:@4410.4]
  assign Multiplexer_Hw_10_io_0 = io_7; // @[Dedicated_PE.scala 121:15:@4409.4]
  assign Multiplexer_Hw_11_io_4 = config_registers_6[13:12]; // @[Dedicated_PE.scala 130:45:@4512.4]
  assign Multiplexer_Hw_11_io_2 = io_15; // @[Dedicated_PE.scala 121:15:@4415.4]
  assign Multiplexer_Hw_11_io_1 = io_11; // @[Dedicated_PE.scala 121:15:@4414.4]
  assign Multiplexer_Hw_11_io_0 = io_7; // @[Dedicated_PE.scala 121:15:@4413.4]
  assign Multiplexer_Hw_12_io_4 = config_registers_6[15:14]; // @[Dedicated_PE.scala 130:45:@4514.4]
  assign Multiplexer_Hw_12_io_2 = io_16; // @[Dedicated_PE.scala 121:15:@4419.4]
  assign Multiplexer_Hw_12_io_1 = io_12; // @[Dedicated_PE.scala 121:15:@4418.4]
  assign Multiplexer_Hw_12_io_0 = io_8; // @[Dedicated_PE.scala 121:15:@4417.4]
  assign Multiplexer_Hw_13_io_4 = config_registers_7[1:0]; // @[Dedicated_PE.scala 130:45:@4516.4]
  assign Multiplexer_Hw_13_io_2 = io_16; // @[Dedicated_PE.scala 121:15:@4423.4]
  assign Multiplexer_Hw_13_io_1 = io_12; // @[Dedicated_PE.scala 121:15:@4422.4]
  assign Multiplexer_Hw_13_io_0 = io_8; // @[Dedicated_PE.scala 121:15:@4421.4]
  assign Multiplexer_Hw_14_io_4 = config_registers_7[3:2]; // @[Dedicated_PE.scala 130:45:@4518.4]
  assign Multiplexer_Hw_14_io_2 = io_16; // @[Dedicated_PE.scala 121:15:@4427.4]
  assign Multiplexer_Hw_14_io_1 = io_12; // @[Dedicated_PE.scala 121:15:@4426.4]
  assign Multiplexer_Hw_14_io_0 = io_8; // @[Dedicated_PE.scala 121:15:@4425.4]
  assign Multiplexer_Hw_15_io_4 = config_registers_7[5:4]; // @[Dedicated_PE.scala 130:45:@4520.4]
  assign Multiplexer_Hw_15_io_2 = io_17; // @[Dedicated_PE.scala 121:15:@4431.4]
  assign Multiplexer_Hw_15_io_1 = io_13; // @[Dedicated_PE.scala 121:15:@4430.4]
  assign Multiplexer_Hw_15_io_0 = io_9; // @[Dedicated_PE.scala 121:15:@4429.4]
  assign Multiplexer_Hw_16_io_4 = config_registers_7[7:6]; // @[Dedicated_PE.scala 130:45:@4522.4]
  assign Multiplexer_Hw_16_io_2 = io_17; // @[Dedicated_PE.scala 121:15:@4435.4]
  assign Multiplexer_Hw_16_io_1 = io_13; // @[Dedicated_PE.scala 121:15:@4434.4]
  assign Multiplexer_Hw_16_io_0 = io_9; // @[Dedicated_PE.scala 121:15:@4433.4]
  assign Multiplexer_Hw_17_io_4 = config_registers_7[9:8]; // @[Dedicated_PE.scala 130:45:@4524.4]
  assign Multiplexer_Hw_17_io_2 = io_17; // @[Dedicated_PE.scala 121:15:@4439.4]
  assign Multiplexer_Hw_17_io_1 = io_13; // @[Dedicated_PE.scala 121:15:@4438.4]
  assign Multiplexer_Hw_17_io_0 = io_9; // @[Dedicated_PE.scala 121:15:@4437.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  config_registers_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  config_registers_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  config_registers_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  config_registers_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  config_registers_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  config_registers_5 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  config_registers_6 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  config_registers_7 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (io_24_write_req) begin
      if (3'h0 == _T_167) begin
        config_registers_0 <= io_24_write_data;
      end
    end
    if (io_24_write_req) begin
      if (3'h1 == _T_167) begin
        config_registers_1 <= io_24_write_data;
      end
    end
    if (io_24_write_req) begin
      if (3'h2 == _T_167) begin
        config_registers_2 <= io_24_write_data;
      end
    end
    if (io_24_write_req) begin
      if (3'h3 == _T_167) begin
        config_registers_3 <= io_24_write_data;
      end
    end
    if (io_24_write_req) begin
      if (3'h4 == _T_167) begin
        config_registers_4 <= io_24_write_data;
      end
    end
    if (io_24_write_req) begin
      if (3'h5 == _T_167) begin
        config_registers_5 <= io_24_write_data;
      end
    end
    if (io_24_write_req) begin
      if (3'h6 == _T_167) begin
        config_registers_6 <= io_24_write_data;
      end
    end
    if (io_24_write_req) begin
      if (3'h7 == _T_167) begin
        config_registers_7 <= io_24_write_data;
      end
    end
  end
endmodule
